//    Xilinx Proprietary Primitive Cell X_UPAD for Verilog
//
// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/xec_libs/data/simprims/X_UPAD.v,v 1.2 2008/10/02 19:01:56 vandanad Exp $
//

`celldefine
`timescale 1 ps/1 ps

module X_UPAD (PAD);

  input PAD;
  parameter LOC = "UNPLACED";
endmodule
