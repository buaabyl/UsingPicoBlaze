///////////////////////////////////////////////////////////
//  Copyright (c) 1995/2006 Xilinx Inc.
//  All Right Reserved.
///////////////////////////////////////////////////////////
//
//   ____   ___
//  /   /\/   / 
// /___/  \  /    Vendor      : Xilinx 
// \  \    \/     Version     : 10.1i
//  \  \          Description : 
//  /  /                      
// /__/   /\      Filename    : X_GTX_DUAL.v
// \  \  /  \     Timestamp   : Tues Nov 13 10:05:08 2007
//  \__\/\__ \                    
//                                 
//  Revision:
//  11/13/07 - Initial version.
//////////////////////////////////////////////////////////////////////////////////

`timescale 1 ps / 1 ps 

module X_GTX_DUAL (
    DFECLKDLYADJMONITOR0,
    DFECLKDLYADJMONITOR1,
    DFEEYEDACMONITOR0,
    DFEEYEDACMONITOR1,
    DFESENSCAL0,
    DFESENSCAL1,
    DFETAP1MONITOR0,
    DFETAP1MONITOR1,
    DFETAP2MONITOR0,
    DFETAP2MONITOR1,
    DFETAP3MONITOR0,
    DFETAP3MONITOR1,
    DFETAP4MONITOR0,
    DFETAP4MONITOR1,
    DO,
    DRDY,
    PHYSTATUS0,
    PHYSTATUS1,
    PLLLKDET,
    REFCLKOUT,
    RESETDONE0,
    RESETDONE1,
    RXBUFSTATUS0,
    RXBUFSTATUS1,
    RXBYTEISALIGNED0,
    RXBYTEISALIGNED1,
    RXBYTEREALIGN0,
    RXBYTEREALIGN1,
    RXCHANBONDSEQ0,
    RXCHANBONDSEQ1,
    RXCHANISALIGNED0,
    RXCHANISALIGNED1,
    RXCHANREALIGN0,
    RXCHANREALIGN1,
    RXCHARISCOMMA0,
    RXCHARISCOMMA1,
    RXCHARISK0,
    RXCHARISK1,
    RXCHBONDO0,
    RXCHBONDO1,
    RXCLKCORCNT0,
    RXCLKCORCNT1,
    RXCOMMADET0,
    RXCOMMADET1,
    RXDATA0,
    RXDATA1,
    RXDATAVALID0,
    RXDATAVALID1,
    RXDISPERR0,
    RXDISPERR1,
    RXELECIDLE0,
    RXELECIDLE1,
    RXHEADER0,
    RXHEADER1,
    RXHEADERVALID0,
    RXHEADERVALID1,
    RXLOSSOFSYNC0,
    RXLOSSOFSYNC1,
    RXNOTINTABLE0,
    RXNOTINTABLE1,
    RXOVERSAMPLEERR0,
    RXOVERSAMPLEERR1,
    RXPRBSERR0,
    RXPRBSERR1,
    RXRECCLK0,
    RXRECCLK1,
    RXRUNDISP0,
    RXRUNDISP1,
    RXSTARTOFSEQ0,
    RXSTARTOFSEQ1,
    RXSTATUS0,
    RXSTATUS1,
    RXVALID0,
    RXVALID1,
    TXBUFSTATUS0,
    TXBUFSTATUS1,
    TXGEARBOXREADY0,
    TXGEARBOXREADY1,
    TXKERR0,
    TXKERR1,
    TXN0,
    TXN1,
    TXOUTCLK0,
    TXOUTCLK1,
    TXP0,
    TXP1,
    TXRUNDISP0,
    TXRUNDISP1,

    CLKIN,
    DADDR,
    DCLK,
    DEN,
    DFECLKDLYADJ0,
    DFECLKDLYADJ1,
    DFETAP10,
    DFETAP11,
    DFETAP20,
    DFETAP21,
    DFETAP30,
    DFETAP31,
    DFETAP40,
    DFETAP41,
    DI,
    DWE,
    GTXRESET,
    GTXTEST,
    INTDATAWIDTH,
    LOOPBACK0,
    LOOPBACK1,
    PLLLKDETEN,
    PLLPOWERDOWN,
    PRBSCNTRESET0,
    PRBSCNTRESET1,
    REFCLKPWRDNB,
    RXBUFRESET0,
    RXBUFRESET1,
    RXCDRRESET0,
    RXCDRRESET1,
    RXCHBONDI0,
    RXCHBONDI1,
    RXCOMMADETUSE0,
    RXCOMMADETUSE1,
    RXDATAWIDTH0,
    RXDATAWIDTH1,
    RXDEC8B10BUSE0,
    RXDEC8B10BUSE1,
    RXENCHANSYNC0,
    RXENCHANSYNC1,
    RXENEQB0,
    RXENEQB1,
    RXENMCOMMAALIGN0,
    RXENMCOMMAALIGN1,
    RXENPCOMMAALIGN0,
    RXENPCOMMAALIGN1,
    RXENPMAPHASEALIGN0,
    RXENPMAPHASEALIGN1,
    RXENPRBSTST0,
    RXENPRBSTST1,
    RXENSAMPLEALIGN0,
    RXENSAMPLEALIGN1,
    RXEQMIX0,
    RXEQMIX1,
    RXEQPOLE0,
    RXEQPOLE1,
    RXGEARBOXSLIP0,
    RXGEARBOXSLIP1,
    RXN0,
    RXN1,
    RXP0,
    RXP1,
    RXPMASETPHASE0,
    RXPMASETPHASE1,
    RXPOLARITY0,
    RXPOLARITY1,
    RXPOWERDOWN0,
    RXPOWERDOWN1,
    RXRESET0,
    RXRESET1,
    RXSLIDE0,
    RXSLIDE1,
    RXUSRCLK0,
    RXUSRCLK1,
    RXUSRCLK20,
    RXUSRCLK21,
    TXBUFDIFFCTRL0,
    TXBUFDIFFCTRL1,
    TXBYPASS8B10B0,
    TXBYPASS8B10B1,
    TXCHARDISPMODE0,
    TXCHARDISPMODE1,
    TXCHARDISPVAL0,
    TXCHARDISPVAL1,
    TXCHARISK0,
    TXCHARISK1,
    TXCOMSTART0,
    TXCOMSTART1,
    TXCOMTYPE0,
    TXCOMTYPE1,
    TXDATA0,
    TXDATA1,
    TXDATAWIDTH0,
    TXDATAWIDTH1,
    TXDETECTRX0,
    TXDETECTRX1,
    TXDIFFCTRL0,
    TXDIFFCTRL1,
    TXELECIDLE0,
    TXELECIDLE1,
    TXENC8B10BUSE0,
    TXENC8B10BUSE1,
    TXENPMAPHASEALIGN0,
    TXENPMAPHASEALIGN1,
    TXENPRBSTST0,
    TXENPRBSTST1,
    TXHEADER0,
    TXHEADER1,
    TXINHIBIT0,
    TXINHIBIT1,
    TXPMASETPHASE0,
    TXPMASETPHASE1,
    TXPOLARITY0,
    TXPOLARITY1,
    TXPOWERDOWN0,
    TXPOWERDOWN1,
    TXPREEMPHASIS0,
    TXPREEMPHASIS1,
    TXRESET0,
    TXRESET1,
    TXSEQUENCE0,
    TXSEQUENCE1,
    TXSTARTSEQ0,
    TXSTARTSEQ1,
    TXUSRCLK0,
    TXUSRCLK1,
    TXUSRCLK20,
    TXUSRCLK21

);


parameter AC_CAP_DIS_0 = "TRUE";
parameter AC_CAP_DIS_1 = "TRUE";
parameter CHAN_BOND_KEEP_ALIGN_0 = "FALSE";
parameter CHAN_BOND_KEEP_ALIGN_1 = "FALSE";
parameter CHAN_BOND_MODE_0 = "OFF";
parameter CHAN_BOND_MODE_1 = "OFF";
parameter CHAN_BOND_SEQ_2_USE_0 = "TRUE";
parameter CHAN_BOND_SEQ_2_USE_1 = "TRUE";
parameter CLKINDC_B = "TRUE";
parameter CLKRCV_TRST = "FALSE";
parameter CLK_CORRECT_USE_0 = "TRUE";
parameter CLK_CORRECT_USE_1 = "TRUE";
parameter CLK_COR_INSERT_IDLE_FLAG_0 = "FALSE";
parameter CLK_COR_INSERT_IDLE_FLAG_1 = "FALSE";
parameter CLK_COR_KEEP_IDLE_0 = "FALSE";
parameter CLK_COR_KEEP_IDLE_1 = "FALSE";
parameter CLK_COR_PRECEDENCE_0 = "TRUE";
parameter CLK_COR_PRECEDENCE_1 = "TRUE";
parameter CLK_COR_SEQ_2_USE_0 = "FALSE";
parameter CLK_COR_SEQ_2_USE_1 = "FALSE";
parameter COMMA_DOUBLE_0 = "FALSE";
parameter COMMA_DOUBLE_1 = "FALSE";
parameter DEC_MCOMMA_DETECT_0 = "TRUE";
parameter DEC_MCOMMA_DETECT_1 = "TRUE";
parameter DEC_PCOMMA_DETECT_0 = "TRUE";
parameter DEC_PCOMMA_DETECT_1 = "TRUE";
parameter DEC_VALID_COMMA_ONLY_0 = "TRUE";
parameter DEC_VALID_COMMA_ONLY_1 = "TRUE";
parameter MCOMMA_DETECT_0 = "TRUE";
parameter MCOMMA_DETECT_1 = "TRUE";
parameter OVERSAMPLE_MODE = "FALSE";
parameter PCI_EXPRESS_MODE_0 = "TRUE";
parameter PCI_EXPRESS_MODE_1 = "TRUE";
parameter PCOMMA_DETECT_0 = "TRUE";
parameter PCOMMA_DETECT_1 = "TRUE";
parameter PLL_FB_DCCEN = "FALSE";
parameter PLL_SATA_0 = "FALSE";
parameter PLL_SATA_1 = "FALSE";
parameter RCV_TERM_GND_0 = "TRUE";
parameter RCV_TERM_GND_1 = "TRUE";
parameter RCV_TERM_VTTRX_0 = "FALSE";
parameter RCV_TERM_VTTRX_1 = "FALSE";
parameter RXGEARBOX_USE_0 = "FALSE";
parameter RXGEARBOX_USE_1 = "FALSE";
parameter RX_BUFFER_USE_0 = "TRUE";
parameter RX_BUFFER_USE_1 = "TRUE";
parameter RX_DECODE_SEQ_MATCH_0 = "TRUE";
parameter RX_DECODE_SEQ_MATCH_1 = "TRUE";
parameter RX_EN_IDLE_HOLD_CDR = "FALSE";
parameter RX_EN_IDLE_HOLD_DFE_0 = "TRUE";
parameter RX_EN_IDLE_HOLD_DFE_1 = "TRUE";
parameter RX_EN_IDLE_RESET_BUF_0 = "TRUE";
parameter RX_EN_IDLE_RESET_BUF_1 = "TRUE";
parameter RX_EN_IDLE_RESET_FR = "TRUE";
parameter RX_EN_IDLE_RESET_PH = "TRUE";
parameter RX_LOSS_OF_SYNC_FSM_0 = "FALSE";
parameter RX_LOSS_OF_SYNC_FSM_1 = "FALSE";
parameter RX_SLIDE_MODE_0 = "PCS";
parameter RX_SLIDE_MODE_1 = "PCS";
parameter RX_STATUS_FMT_0 = "PCIE";
parameter RX_STATUS_FMT_1 = "PCIE";
parameter RX_XCLK_SEL_0 = "RXREC";
parameter RX_XCLK_SEL_1 = "RXREC";
parameter SIM_PLL_PERDIV2 = 9'h190;
parameter SIM_RECEIVER_DETECT_PASS_0 = "FALSE";
parameter SIM_RECEIVER_DETECT_PASS_1 = "FALSE";
parameter TERMINATION_OVRD = "FALSE";
parameter TXGEARBOX_USE_0 = "FALSE";
parameter TXGEARBOX_USE_1 = "FALSE";
parameter TX_BUFFER_USE_0 = "TRUE";
parameter TX_BUFFER_USE_1 = "TRUE";
parameter TX_XCLK_SEL_0 = "TXUSR";
parameter TX_XCLK_SEL_1 = "TXUSR";
parameter [11:0] TRANS_TIME_FROM_P2_0 = 12'h03c;
parameter [11:0] TRANS_TIME_FROM_P2_1 = 12'h03c;
parameter [13:0] TX_DETECT_RX_CFG_0 = 14'h1832;
parameter [13:0] TX_DETECT_RX_CFG_1 = 14'h1832;
parameter [19:0] PMA_TX_CFG_0 = 20'h00082;
parameter [19:0] PMA_TX_CFG_1 = 20'h00082;
parameter [1:0] CM_TRIM_0 = 2'b10;
parameter [1:0] CM_TRIM_1 = 2'b10;
parameter [23:0] PLL_COM_CFG = 24'h21680a;
parameter [24:0] PMA_RX_CFG_0 = 25'h05ce109;
parameter [24:0] PMA_RX_CFG_1 = 25'h05ce109;
parameter [26:0] PMA_CDR_SCAN_0 = 27'h6c08040;
parameter [26:0] PMA_CDR_SCAN_1 = 27'h6c08040;
parameter [2:0] GEARBOX_ENDEC_0 = 3'b000;
parameter [2:0] GEARBOX_ENDEC_1 = 3'b000;
parameter [2:0] OOBDETECT_THRESHOLD_0 = 3'b111;
parameter [2:0] OOBDETECT_THRESHOLD_1 = 3'b111;
parameter [2:0] PLL_LKDET_CFG = 3'b111;
parameter [2:0] PLL_TDCC_CFG = 3'b000;
parameter [2:0] SATA_BURST_VAL_0 = 3'b100;
parameter [2:0] SATA_BURST_VAL_1 = 3'b100;
parameter [2:0] SATA_IDLE_VAL_0 = 3'b011;
parameter [2:0] SATA_IDLE_VAL_1 = 3'b011;
parameter [2:0] TXRX_INVERT_0 = 3'b000;
parameter [2:0] TXRX_INVERT_1 = 3'b000;
parameter [2:0] TX_IDLE_DELAY_0 = 3'b010;
parameter [2:0] TX_IDLE_DELAY_1 = 3'b010;
parameter [31:0] PRBS_ERR_THRESHOLD_0 = 32'h1;
parameter [31:0] PRBS_ERR_THRESHOLD_1 = 32'h1;
parameter [3:0] CHAN_BOND_SEQ_1_ENABLE_0 = 4'b1111;
parameter [3:0] CHAN_BOND_SEQ_1_ENABLE_1 = 4'b1111;
parameter [3:0] CHAN_BOND_SEQ_2_ENABLE_0 = 4'b1111;
parameter [3:0] CHAN_BOND_SEQ_2_ENABLE_1 = 4'b1111;
parameter [3:0] CLK_COR_SEQ_1_ENABLE_0 = 4'b1111;
parameter [3:0] CLK_COR_SEQ_1_ENABLE_1 = 4'b1111;
parameter [3:0] CLK_COR_SEQ_2_ENABLE_0 = 4'b1111;
parameter [3:0] CLK_COR_SEQ_2_ENABLE_1 = 4'b1111;
parameter [3:0] COM_BURST_VAL_0 = 4'b1111;
parameter [3:0] COM_BURST_VAL_1 = 4'b1111;
parameter [3:0] RX_IDLE_HI_CNT_0 = 4'b1000;
parameter [3:0] RX_IDLE_HI_CNT_1 = 4'b1000;
parameter [3:0] RX_IDLE_LO_CNT_0 = 4'b0000;
parameter [3:0] RX_IDLE_LO_CNT_1 = 4'b0000;
parameter [4:0] CDR_PH_ADJ_TIME = 5'b01010;
parameter [4:0] DFE_CAL_TIME = 5'b00110;
parameter [4:0] TERMINATION_CTRL = 5'b10100;
parameter [68:0] PMA_COM_CFG = 69'h0;
parameter [6:0] PMA_RXSYNC_CFG_0 = 7'h0;
parameter [6:0] PMA_RXSYNC_CFG_1 = 7'h0;
parameter [7:0] PLL_CP_CFG = 8'h00;
parameter [7:0] TRANS_TIME_NON_P2_0 = 8'h19;
parameter [7:0] TRANS_TIME_NON_P2_1 = 8'h19;
parameter [9:0] CHAN_BOND_SEQ_1_1_0 = 10'b0001001010;
parameter [9:0] CHAN_BOND_SEQ_1_1_1 = 10'b0001001010;
parameter [9:0] CHAN_BOND_SEQ_1_2_0 = 10'b0001001010;
parameter [9:0] CHAN_BOND_SEQ_1_2_1 = 10'b0001001010;
parameter [9:0] CHAN_BOND_SEQ_1_3_0 = 10'b0001001010;
parameter [9:0] CHAN_BOND_SEQ_1_3_1 = 10'b0001001010;
parameter [9:0] CHAN_BOND_SEQ_1_4_0 = 10'b0110111100;
parameter [9:0] CHAN_BOND_SEQ_1_4_1 = 10'b0110111100;
parameter [9:0] CHAN_BOND_SEQ_2_1_0 = 10'b0110111100;
parameter [9:0] CHAN_BOND_SEQ_2_1_1 = 10'b0110111100;
parameter [9:0] CHAN_BOND_SEQ_2_2_0 = 10'b0100111100;
parameter [9:0] CHAN_BOND_SEQ_2_2_1 = 10'b0100111100;
parameter [9:0] CHAN_BOND_SEQ_2_3_0 = 10'b0100111100;
parameter [9:0] CHAN_BOND_SEQ_2_3_1 = 10'b0100111100;
parameter [9:0] CHAN_BOND_SEQ_2_4_0 = 10'b0100111100;
parameter [9:0] CHAN_BOND_SEQ_2_4_1 = 10'b0100111100;
parameter [9:0] CLK_COR_SEQ_1_1_0 = 10'b0100011100;
parameter [9:0] CLK_COR_SEQ_1_1_1 = 10'b0100011100;
parameter [9:0] CLK_COR_SEQ_1_2_0 = 10'b0;
parameter [9:0] CLK_COR_SEQ_1_2_1 = 10'b0;
parameter [9:0] CLK_COR_SEQ_1_3_0 = 10'b0;
parameter [9:0] CLK_COR_SEQ_1_3_1 = 10'b0;
parameter [9:0] CLK_COR_SEQ_1_4_0 = 10'b0;
parameter [9:0] CLK_COR_SEQ_1_4_1 = 10'b0;
parameter [9:0] CLK_COR_SEQ_2_1_0 = 10'b0;
parameter [9:0] CLK_COR_SEQ_2_1_1 = 10'b0;
parameter [9:0] CLK_COR_SEQ_2_2_0 = 10'b0;
parameter [9:0] CLK_COR_SEQ_2_2_1 = 10'b0;
parameter [9:0] CLK_COR_SEQ_2_3_0 = 10'b0;
parameter [9:0] CLK_COR_SEQ_2_3_1 = 10'b0;
parameter [9:0] CLK_COR_SEQ_2_4_0 = 10'b0;
parameter [9:0] CLK_COR_SEQ_2_4_1 = 10'b0;
parameter [9:0] COMMA_10B_ENABLE_0 = 10'b1111111111;
parameter [9:0] COMMA_10B_ENABLE_1 = 10'b1111111111;
parameter [9:0] DFE_CFG_0 = 10'b0001111011;
parameter [9:0] DFE_CFG_1 = 10'b0001111011;
parameter [9:0] MCOMMA_10B_VALUE_0 = 10'b1010000011;
parameter [9:0] MCOMMA_10B_VALUE_1 = 10'b1010000011;
parameter [9:0] PCOMMA_10B_VALUE_0 = 10'b0101111100;
parameter [9:0] PCOMMA_10B_VALUE_1 = 10'b0101111100;
parameter [9:0] TRANS_TIME_TO_P2_0 = 10'h064;
parameter [9:0] TRANS_TIME_TO_P2_1 = 10'h064;
parameter  ALIGN_COMMA_WORD_0 = 1;
parameter  ALIGN_COMMA_WORD_1 = 1;
parameter  CB2_INH_CC_PERIOD_0 = 8;
parameter  CB2_INH_CC_PERIOD_1 = 8;
parameter  CHAN_BOND_1_MAX_SKEW_0 = 7;
parameter  CHAN_BOND_1_MAX_SKEW_1 = 7;
parameter  CHAN_BOND_2_MAX_SKEW_0 = 1;
parameter  CHAN_BOND_2_MAX_SKEW_1 = 1;
parameter  CHAN_BOND_LEVEL_0 = 0;
parameter  CHAN_BOND_LEVEL_1 = 0;
parameter  CHAN_BOND_SEQ_LEN_0 = 4;
parameter  CHAN_BOND_SEQ_LEN_1 = 4;
parameter  CLK25_DIVIDER = 4;
parameter  CLK_COR_ADJ_LEN_0 = 1;
parameter  CLK_COR_ADJ_LEN_1 = 1;
parameter  CLK_COR_DET_LEN_0 = 1;
parameter  CLK_COR_DET_LEN_1 = 1;
parameter  CLK_COR_MAX_LAT_0 = 18;
parameter  CLK_COR_MAX_LAT_1 = 18;
parameter  CLK_COR_MIN_LAT_0 = 16;
parameter  CLK_COR_MIN_LAT_1 = 16;
parameter  CLK_COR_REPEAT_WAIT_0 = 5;
parameter  CLK_COR_REPEAT_WAIT_1 = 5;
parameter  OOB_CLK_DIVIDER = 4;
parameter  PLL_DIVSEL_FB = 5;
parameter  PLL_DIVSEL_REF = 2;
parameter  PLL_RXDIVSEL_OUT_0 = 1;
parameter  PLL_RXDIVSEL_OUT_1 = 1;
parameter  PLL_TXDIVSEL_OUT_0 = 1;
parameter  PLL_TXDIVSEL_OUT_1 = 1;
parameter  RX_LOS_INVALID_INCR_0 = 8;
parameter  RX_LOS_INVALID_INCR_1 = 8;
parameter  RX_LOS_THRESHOLD_0 = 128;
parameter  RX_LOS_THRESHOLD_1 = 128;
parameter  SATA_MAX_BURST_0 = 7;
parameter  SATA_MAX_BURST_1 = 7;
parameter  SATA_MAX_INIT_0 = 22;
parameter  SATA_MAX_INIT_1 = 22;
parameter  SATA_MAX_WAKE_0 = 7;
parameter  SATA_MAX_WAKE_1 = 7;
parameter  SATA_MIN_BURST_0 = 4;
parameter  SATA_MIN_BURST_1 = 4;
parameter  SATA_MIN_INIT_0 = 12;
parameter  SATA_MIN_INIT_1 = 12;
parameter  SATA_MIN_WAKE_0 = 4;
parameter  SATA_MIN_WAKE_1 = 4;
parameter  SIM_GTXRESET_SPEEDUP = 0;
parameter  TERMINATION_IMP_0 = 50;
parameter  TERMINATION_IMP_1 = 50;
parameter LOC = "UNPLACED";
localparam in_delay =  0;
localparam out_delay = 0;
localparam CLK_DELAY = 0;

output DRDY;
output PHYSTATUS0;
output PHYSTATUS1;
output PLLLKDET;
output REFCLKOUT;
output RESETDONE0;
output RESETDONE1;
output RXBYTEISALIGNED0;
output RXBYTEISALIGNED1;
output RXBYTEREALIGN0;
output RXBYTEREALIGN1;
output RXCHANBONDSEQ0;
output RXCHANBONDSEQ1;
output RXCHANISALIGNED0;
output RXCHANISALIGNED1;
output RXCHANREALIGN0;
output RXCHANREALIGN1;
output RXCOMMADET0;
output RXCOMMADET1;
output RXDATAVALID0;
output RXDATAVALID1;
output RXELECIDLE0;
output RXELECIDLE1;
output RXHEADERVALID0;
output RXHEADERVALID1;
output RXOVERSAMPLEERR0;
output RXOVERSAMPLEERR1;
output RXPRBSERR0;
output RXPRBSERR1;
output RXRECCLK0;
output RXRECCLK1;
output RXSTARTOFSEQ0;
output RXSTARTOFSEQ1;
output RXVALID0;
output RXVALID1;
output TXGEARBOXREADY0;
output TXGEARBOXREADY1;
output TXN0;
output TXN1;
output TXOUTCLK0;
output TXOUTCLK1;
output TXP0;
output TXP1;
output [15:0] DO;
output [1:0] RXLOSSOFSYNC0;
output [1:0] RXLOSSOFSYNC1;
output [1:0] TXBUFSTATUS0;
output [1:0] TXBUFSTATUS1;
output [2:0] DFESENSCAL0;
output [2:0] DFESENSCAL1;
output [2:0] RXBUFSTATUS0;
output [2:0] RXBUFSTATUS1;
output [2:0] RXCLKCORCNT0;
output [2:0] RXCLKCORCNT1;
output [2:0] RXHEADER0;
output [2:0] RXHEADER1;
output [2:0] RXSTATUS0;
output [2:0] RXSTATUS1;
output [31:0] RXDATA0;
output [31:0] RXDATA1;
output [3:0] DFETAP3MONITOR0;
output [3:0] DFETAP3MONITOR1;
output [3:0] DFETAP4MONITOR0;
output [3:0] DFETAP4MONITOR1;
output [3:0] RXCHARISCOMMA0;
output [3:0] RXCHARISCOMMA1;
output [3:0] RXCHARISK0;
output [3:0] RXCHARISK1;
output [3:0] RXCHBONDO0;
output [3:0] RXCHBONDO1;
output [3:0] RXDISPERR0;
output [3:0] RXDISPERR1;
output [3:0] RXNOTINTABLE0;
output [3:0] RXNOTINTABLE1;
output [3:0] RXRUNDISP0;
output [3:0] RXRUNDISP1;
output [3:0] TXKERR0;
output [3:0] TXKERR1;
output [3:0] TXRUNDISP0;
output [3:0] TXRUNDISP1;
output [4:0] DFEEYEDACMONITOR0;
output [4:0] DFEEYEDACMONITOR1;
output [4:0] DFETAP1MONITOR0;
output [4:0] DFETAP1MONITOR1;
output [4:0] DFETAP2MONITOR0;
output [4:0] DFETAP2MONITOR1;
output [5:0] DFECLKDLYADJMONITOR0;
output [5:0] DFECLKDLYADJMONITOR1;

input CLKIN;
input DCLK;
input DEN;
input DWE;
input GTXRESET;
input INTDATAWIDTH;
input PLLLKDETEN;
input PLLPOWERDOWN;
input PRBSCNTRESET0;
input PRBSCNTRESET1;
input REFCLKPWRDNB;
input RXBUFRESET0;
input RXBUFRESET1;
input RXCDRRESET0;
input RXCDRRESET1;
input RXCOMMADETUSE0;
input RXCOMMADETUSE1;
input RXDEC8B10BUSE0;
input RXDEC8B10BUSE1;
input RXENCHANSYNC0;
input RXENCHANSYNC1;
input RXENEQB0;
input RXENEQB1;
input RXENMCOMMAALIGN0;
input RXENMCOMMAALIGN1;
input RXENPCOMMAALIGN0;
input RXENPCOMMAALIGN1;
input RXENPMAPHASEALIGN0;
input RXENPMAPHASEALIGN1;
input RXENSAMPLEALIGN0;
input RXENSAMPLEALIGN1;
input RXGEARBOXSLIP0;
input RXGEARBOXSLIP1;
input RXN0;
input RXN1;
input RXP0;
input RXP1;
input RXPMASETPHASE0;
input RXPMASETPHASE1;
input RXPOLARITY0;
input RXPOLARITY1;
input RXRESET0;
input RXRESET1;
input RXSLIDE0;
input RXSLIDE1;
input RXUSRCLK0;
input RXUSRCLK1;
input RXUSRCLK20;
input RXUSRCLK21;
input TXCOMSTART0;
input TXCOMSTART1;
input TXCOMTYPE0;
input TXCOMTYPE1;
input TXDETECTRX0;
input TXDETECTRX1;
input TXELECIDLE0;
input TXELECIDLE1;
input TXENC8B10BUSE0;
input TXENC8B10BUSE1;
input TXENPMAPHASEALIGN0;
input TXENPMAPHASEALIGN1;
input TXINHIBIT0;
input TXINHIBIT1;
input TXPMASETPHASE0;
input TXPMASETPHASE1;
input TXPOLARITY0;
input TXPOLARITY1;
input TXRESET0;
input TXRESET1;
input TXSTARTSEQ0;
input TXSTARTSEQ1;
input TXUSRCLK0;
input TXUSRCLK1;
input TXUSRCLK20;
input TXUSRCLK21;
input [13:0] GTXTEST;
input [15:0] DI;
input [1:0] RXDATAWIDTH0;
input [1:0] RXDATAWIDTH1;
input [1:0] RXENPRBSTST0;
input [1:0] RXENPRBSTST1;
input [1:0] RXEQMIX0;
input [1:0] RXEQMIX1;
input [1:0] RXPOWERDOWN0;
input [1:0] RXPOWERDOWN1;
input [1:0] TXDATAWIDTH0;
input [1:0] TXDATAWIDTH1;
input [1:0] TXENPRBSTST0;
input [1:0] TXENPRBSTST1;
input [1:0] TXPOWERDOWN0;
input [1:0] TXPOWERDOWN1;
input [2:0] LOOPBACK0;
input [2:0] LOOPBACK1;
input [2:0] TXBUFDIFFCTRL0;
input [2:0] TXBUFDIFFCTRL1;
input [2:0] TXDIFFCTRL0;
input [2:0] TXDIFFCTRL1;
input [2:0] TXHEADER0;
input [2:0] TXHEADER1;
input [31:0] TXDATA0;
input [31:0] TXDATA1;
input [3:0] DFETAP30;
input [3:0] DFETAP31;
input [3:0] DFETAP40;
input [3:0] DFETAP41;
input [3:0] RXCHBONDI0;
input [3:0] RXCHBONDI1;
input [3:0] RXEQPOLE0;
input [3:0] RXEQPOLE1;
input [3:0] TXBYPASS8B10B0;
input [3:0] TXBYPASS8B10B1;
input [3:0] TXCHARDISPMODE0;
input [3:0] TXCHARDISPMODE1;
input [3:0] TXCHARDISPVAL0;
input [3:0] TXCHARDISPVAL1;
input [3:0] TXCHARISK0;
input [3:0] TXCHARISK1;
input [3:0] TXPREEMPHASIS0;
input [3:0] TXPREEMPHASIS1;
input [4:0] DFETAP10;
input [4:0] DFETAP11;
input [4:0] DFETAP20;
input [4:0] DFETAP21;
input [5:0] DFECLKDLYADJ0;
input [5:0] DFECLKDLYADJ1;
input [6:0] DADDR;
input [6:0] TXSEQUENCE0;
input [6:0] TXSEQUENCE1;

endmodule
