///////////////////////////////////////////////////////////
//  Copyright (c) 1995/2006 Xilinx Inc.
//  All Right Reserved.
///////////////////////////////////////////////////////////
//
//   ____   ___
//  /   /\/   / 
// /___/  \  /    Vendor      : Xilinx 
// \  \    \/     Version : 10.1
//  \  \          Description : Xilinx Formal Library Component
//  /  /                        PCI Express
// /__/   /\      Filename    : PCIE_INTERNAL_1_1.v
// \  \  /  \     Timestamp   : Mon Nov 12 2007   
//  \__\/\__ \                    
//                                 
//  Revision:
//    11/12/07 - Initial version.
///////////////////////////////////////////////////////////

`timescale 1 ps / 1 ps 

module PCIE_INTERNAL_1_1 (
    BUSMASTERENABLE,
    CRMDOHOTRESETN,
    CRMPWRSOFTRESETN,
    CRMRXHOTRESETN,
    DLLTXPMDLLPOUTSTANDING,
    INTERRUPTDISABLE,
    IOSPACEENABLE,
    L0ASAUTONOMOUSINITCOMPLETED,
    L0ATTENTIONINDICATORCONTROL,
    L0CFGLOOPBACKACK,
    L0COMPLETERID,
    L0CORRERRMSGRCVD,
    L0DLLASRXSTATE,
    L0DLLASTXSTATE,
    L0DLLERRORVECTOR,
    L0DLLRXACKOUTSTANDING,
    L0DLLTXNONFCOUTSTANDING,
    L0DLLTXOUTSTANDING,
    L0DLLVCSTATUS,
    L0DLUPDOWN,
    L0ERRMSGREQID,
    L0FATALERRMSGRCVD,
    L0FIRSTCFGWRITEOCCURRED,
    L0FWDCORRERROUT,
    L0FWDFATALERROUT,
    L0FWDNONFATALERROUT,
    L0LTSSMSTATE,
    L0MACENTEREDL0,
    L0MACLINKTRAINING,
    L0MACLINKUP,
    L0MACNEGOTIATEDLINKWIDTH,
    L0MACNEWSTATEACK,
    L0MACRXL0SSTATE,
    L0MACUPSTREAMDOWNSTREAM,
    L0MCFOUND,
    L0MSIENABLE0,
    L0MULTIMSGEN0,
    L0NONFATALERRMSGRCVD,
    L0PMEACK,
    L0PMEEN,
    L0PMEREQOUT,
    L0POWERCONTROLLERCONTROL,
    L0POWERINDICATORCONTROL,
    L0PWRINHIBITTRANSFERS,
    L0PWRL1STATE,
    L0PWRL23READYDEVICE,
    L0PWRL23READYSTATE,
    L0PWRSTATE0,
    L0PWRTURNOFFREQ,
    L0PWRTXL0SSTATE,
    L0RECEIVEDASSERTINTALEGACYINT,
    L0RECEIVEDASSERTINTBLEGACYINT,
    L0RECEIVEDASSERTINTCLEGACYINT,
    L0RECEIVEDASSERTINTDLEGACYINT,
    L0RECEIVEDDEASSERTINTALEGACYINT,
    L0RECEIVEDDEASSERTINTBLEGACYINT,
    L0RECEIVEDDEASSERTINTCLEGACYINT,
    L0RECEIVEDDEASSERTINTDLEGACYINT,
    L0RXBEACON,
    L0RXDLLFCCMPLMCCRED,
    L0RXDLLFCCMPLMCUPDATE,
    L0RXDLLFCNPOSTBYPCRED,
    L0RXDLLFCNPOSTBYPUPDATE,
    L0RXDLLFCPOSTORDCRED,
    L0RXDLLFCPOSTORDUPDATE,
    L0RXDLLPM,
    L0RXDLLPMTYPE,
    L0RXDLLSBFCDATA,
    L0RXDLLSBFCUPDATE,
    L0RXDLLTLPECRCOK,
    L0RXDLLTLPEND,
    L0RXMACLINKERROR,
    L0STATSCFGOTHERRECEIVED,
    L0STATSCFGOTHERTRANSMITTED,
    L0STATSCFGRECEIVED,
    L0STATSCFGTRANSMITTED,
    L0STATSDLLPRECEIVED,
    L0STATSDLLPTRANSMITTED,
    L0STATSOSRECEIVED,
    L0STATSOSTRANSMITTED,
    L0STATSTLPRECEIVED,
    L0STATSTLPTRANSMITTED,
    L0TOGGLEELECTROMECHANICALINTERLOCK,
    L0TRANSFORMEDVC,
    L0TXDLLFCCMPLMCUPDATED,
    L0TXDLLFCNPOSTBYPUPDATED,
    L0TXDLLFCPOSTORDUPDATED,
    L0TXDLLPMUPDATED,
    L0TXDLLSBFCUPDATED,
    L0UCBYPFOUND,
    L0UCORDFOUND,
    L0UNLOCKRECEIVED,
    LLKRX4DWHEADERN,
    LLKRXCHCOMPLETIONAVAILABLEN,
    LLKRXCHCOMPLETIONPARTIALN,
    LLKRXCHCONFIGAVAILABLEN,
    LLKRXCHCONFIGPARTIALN,
    LLKRXCHNONPOSTEDAVAILABLEN,
    LLKRXCHNONPOSTEDPARTIALN,
    LLKRXCHPOSTEDAVAILABLEN,
    LLKRXCHPOSTEDPARTIALN,
    LLKRXDATA,
    LLKRXECRCBADN,
    LLKRXEOFN,
    LLKRXEOPN,
    LLKRXPREFERREDTYPE,
    LLKRXSOFN,
    LLKRXSOPN,
    LLKRXSRCDSCN,
    LLKRXSRCLASTREQN,
    LLKRXSRCRDYN,
    LLKRXVALIDN,
    LLKTCSTATUS,
    LLKTXCHANSPACE,
    LLKTXCHCOMPLETIONREADYN,
    LLKTXCHNONPOSTEDREADYN,
    LLKTXCHPOSTEDREADYN,
    LLKTXCONFIGREADYN,
    LLKTXDSTRDYN,
    MAXPAYLOADSIZE,
    MAXREADREQUESTSIZE,
    MEMSPACEENABLE,
    MGMTPSO,
    MGMTRDATA,
    MGMTSTATSCREDIT,
    MIMDLLBRADD,
    MIMDLLBREN,
    MIMDLLBWADD,
    MIMDLLBWDATA,
    MIMDLLBWEN,
    MIMRXBRADD,
    MIMRXBREN,
    MIMRXBWADD,
    MIMRXBWDATA,
    MIMRXBWEN,
    MIMTXBRADD,
    MIMTXBREN,
    MIMTXBWADD,
    MIMTXBWDATA,
    MIMTXBWEN,
    PARITYERRORRESPONSE,
    PIPEDESKEWLANESL0,
    PIPEDESKEWLANESL1,
    PIPEDESKEWLANESL2,
    PIPEDESKEWLANESL3,
    PIPEDESKEWLANESL4,
    PIPEDESKEWLANESL5,
    PIPEDESKEWLANESL6,
    PIPEDESKEWLANESL7,
    PIPEPOWERDOWNL0,
    PIPEPOWERDOWNL1,
    PIPEPOWERDOWNL2,
    PIPEPOWERDOWNL3,
    PIPEPOWERDOWNL4,
    PIPEPOWERDOWNL5,
    PIPEPOWERDOWNL6,
    PIPEPOWERDOWNL7,
    PIPERESETL0,
    PIPERESETL1,
    PIPERESETL2,
    PIPERESETL3,
    PIPERESETL4,
    PIPERESETL5,
    PIPERESETL6,
    PIPERESETL7,
    PIPERXPOLARITYL0,
    PIPERXPOLARITYL1,
    PIPERXPOLARITYL2,
    PIPERXPOLARITYL3,
    PIPERXPOLARITYL4,
    PIPERXPOLARITYL5,
    PIPERXPOLARITYL6,
    PIPERXPOLARITYL7,
    PIPETXCOMPLIANCEL0,
    PIPETXCOMPLIANCEL1,
    PIPETXCOMPLIANCEL2,
    PIPETXCOMPLIANCEL3,
    PIPETXCOMPLIANCEL4,
    PIPETXCOMPLIANCEL5,
    PIPETXCOMPLIANCEL6,
    PIPETXCOMPLIANCEL7,
    PIPETXDATAKL0,
    PIPETXDATAKL1,
    PIPETXDATAKL2,
    PIPETXDATAKL3,
    PIPETXDATAKL4,
    PIPETXDATAKL5,
    PIPETXDATAKL6,
    PIPETXDATAKL7,
    PIPETXDATAL0,
    PIPETXDATAL1,
    PIPETXDATAL2,
    PIPETXDATAL3,
    PIPETXDATAL4,
    PIPETXDATAL5,
    PIPETXDATAL6,
    PIPETXDATAL7,
    PIPETXDETECTRXLOOPBACKL0,
    PIPETXDETECTRXLOOPBACKL1,
    PIPETXDETECTRXLOOPBACKL2,
    PIPETXDETECTRXLOOPBACKL3,
    PIPETXDETECTRXLOOPBACKL4,
    PIPETXDETECTRXLOOPBACKL5,
    PIPETXDETECTRXLOOPBACKL6,
    PIPETXDETECTRXLOOPBACKL7,
    PIPETXELECIDLEL0,
    PIPETXELECIDLEL1,
    PIPETXELECIDLEL2,
    PIPETXELECIDLEL3,
    PIPETXELECIDLEL4,
    PIPETXELECIDLEL5,
    PIPETXELECIDLEL6,
    PIPETXELECIDLEL7,
    SERRENABLE,
    URREPORTINGENABLE,

    AUXPOWER,
    CFGNEGOTIATEDLINKWIDTH,
    COMPLIANCEAVOID,
    CRMCFGBRIDGEHOTRESET,
    CRMCORECLK,
    CRMCORECLKDLO,
    CRMCORECLKRXO,
    CRMCORECLKTXO,
    CRMLINKRSTN,
    CRMMACRSTN,
    CRMMGMTRSTN,
    CRMNVRSTN,
    CRMTXHOTRESETN,
    CRMURSTN,
    CRMUSERCFGRSTN,
    CRMUSERCLK,
    CRMUSERCLKRXO,
    CRMUSERCLKTXO,
    CROSSLINKSEED,
    L0ACKNAKTIMERADJUSTMENT,
    L0ALLDOWNPORTSINL1,
    L0ALLDOWNRXPORTSINL0S,
    L0ASE,
    L0ASPORTCOUNT,
    L0ASTURNPOOLBITSCONSUMED,
    L0ATTENTIONBUTTONPRESSED,
    L0CFGASSPANTREEOWNEDSTATE,
    L0CFGASSTATECHANGECMD,
    L0CFGDISABLESCRAMBLE,
    L0CFGEXTENDEDSYNC,
    L0CFGL0SENTRYENABLE,
    L0CFGL0SENTRYSUP,
    L0CFGL0SEXITLAT,
    L0CFGLINKDISABLE,
    L0CFGLOOPBACKMASTER,
    L0CFGNEGOTIATEDMAXP,
    L0CFGVCENABLE,
    L0CFGVCID,
    L0DLLHOLDLINKUP,
    L0ELECTROMECHANICALINTERLOCKENGAGED,
    L0FWDASSERTINTALEGACYINT,
    L0FWDASSERTINTBLEGACYINT,
    L0FWDASSERTINTCLEGACYINT,
    L0FWDASSERTINTDLEGACYINT,
    L0FWDCORRERRIN,
    L0FWDDEASSERTINTALEGACYINT,
    L0FWDDEASSERTINTBLEGACYINT,
    L0FWDDEASSERTINTCLEGACYINT,
    L0FWDDEASSERTINTDLEGACYINT,
    L0FWDFATALERRIN,
    L0FWDNONFATALERRIN,
    L0LEGACYINTFUNCT0,
    L0MRLSENSORCLOSEDN,
    L0MSIREQUEST0,
    L0PACKETHEADERFROMUSER,
    L0PMEREQIN,
    L0PORTNUMBER,
    L0POWERFAULTDETECTED,
    L0PRESENCEDETECTSLOTEMPTYN,
    L0PWRNEWSTATEREQ,
    L0PWRNEXTLINKSTATE,
    L0REPLAYTIMERADJUSTMENT,
    L0ROOTTURNOFFREQ,
    L0RXTLTLPNONINITIALIZEDVC,
    L0SENDUNLOCKMESSAGE,
    L0SETCOMPLETERABORTERROR,
    L0SETCOMPLETIONTIMEOUTCORRERROR,
    L0SETCOMPLETIONTIMEOUTUNCORRERROR,
    L0SETDETECTEDCORRERROR,
    L0SETDETECTEDFATALERROR,
    L0SETDETECTEDNONFATALERROR,
    L0SETLINKDETECTEDPARITYERROR,
    L0SETLINKMASTERDATAPARITY,
    L0SETLINKRECEIVEDMASTERABORT,
    L0SETLINKRECEIVEDTARGETABORT,
    L0SETLINKSIGNALLEDTARGETABORT,
    L0SETLINKSYSTEMERROR,
    L0SETUNEXPECTEDCOMPLETIONCORRERROR,
    L0SETUNEXPECTEDCOMPLETIONUNCORRERROR,
    L0SETUNSUPPORTEDREQUESTNONPOSTEDERROR,
    L0SETUNSUPPORTEDREQUESTOTHERERROR,
    L0SETUSERDETECTEDPARITYERROR,
    L0SETUSERMASTERDATAPARITY,
    L0SETUSERRECEIVEDMASTERABORT,
    L0SETUSERRECEIVEDTARGETABORT,
    L0SETUSERSIGNALLEDTARGETABORT,
    L0SETUSERSYSTEMERROR,
    L0TLASFCCREDSTARVATION,
    L0TLLINKRETRAIN,
    L0TRANSACTIONSPENDING,
    L0TXBEACON,
    L0TXCFGPM,
    L0TXCFGPMTYPE,
    L0TXTLFCCMPLMCCRED,
    L0TXTLFCCMPLMCUPDATE,
    L0TXTLFCNPOSTBYPCRED,
    L0TXTLFCNPOSTBYPUPDATE,
    L0TXTLFCPOSTORDCRED,
    L0TXTLFCPOSTORDUPDATE,
    L0TXTLSBFCDATA,
    L0TXTLSBFCUPDATE,
    L0TXTLTLPDATA,
    L0TXTLTLPEDB,
    L0TXTLTLPENABLE,
    L0TXTLTLPEND,
    L0TXTLTLPLATENCY,
    L0TXTLTLPREQ,
    L0TXTLTLPREQEND,
    L0TXTLTLPWIDTH,
    L0UPSTREAMRXPORTINL0S,
    L0VC0PREVIEWEXPAND,
    L0WAKEN,
    LLKRXCHFIFO,
    LLKRXCHTC,
    LLKRXDSTCONTREQN,
    LLKRXDSTREQN,
    LLKTX4DWHEADERN,
    LLKTXCHFIFO,
    LLKTXCHTC,
    LLKTXCOMPLETEN,
    LLKTXCREATEECRCN,
    LLKTXDATA,
    LLKTXENABLEN,
    LLKTXEOFN,
    LLKTXEOPN,
    LLKTXSOFN,
    LLKTXSOPN,
    LLKTXSRCDSCN,
    LLKTXSRCRDYN,
    MAINPOWER,
    MGMTADDR,
    MGMTBWREN,
    MGMTRDEN,
    MGMTSTATSCREDITSEL,
    MGMTWDATA,
    MGMTWREN,
    MIMDLLBRDATA,
    MIMRXBRDATA,
    MIMTXBRDATA,
    PIPEPHYSTATUSL0,
    PIPEPHYSTATUSL1,
    PIPEPHYSTATUSL2,
    PIPEPHYSTATUSL3,
    PIPEPHYSTATUSL4,
    PIPEPHYSTATUSL5,
    PIPEPHYSTATUSL6,
    PIPEPHYSTATUSL7,
    PIPERXCHANISALIGNEDL0,
    PIPERXCHANISALIGNEDL1,
    PIPERXCHANISALIGNEDL2,
    PIPERXCHANISALIGNEDL3,
    PIPERXCHANISALIGNEDL4,
    PIPERXCHANISALIGNEDL5,
    PIPERXCHANISALIGNEDL6,
    PIPERXCHANISALIGNEDL7,
    PIPERXDATAKL0,
    PIPERXDATAKL1,
    PIPERXDATAKL2,
    PIPERXDATAKL3,
    PIPERXDATAKL4,
    PIPERXDATAKL5,
    PIPERXDATAKL6,
    PIPERXDATAKL7,
    PIPERXDATAL0,
    PIPERXDATAL1,
    PIPERXDATAL2,
    PIPERXDATAL3,
    PIPERXDATAL4,
    PIPERXDATAL5,
    PIPERXDATAL6,
    PIPERXDATAL7,
    PIPERXELECIDLEL0,
    PIPERXELECIDLEL1,
    PIPERXELECIDLEL2,
    PIPERXELECIDLEL3,
    PIPERXELECIDLEL4,
    PIPERXELECIDLEL5,
    PIPERXELECIDLEL6,
    PIPERXELECIDLEL7,
    PIPERXSTATUSL0,
    PIPERXSTATUSL1,
    PIPERXSTATUSL2,
    PIPERXSTATUSL3,
    PIPERXSTATUSL4,
    PIPERXSTATUSL5,
    PIPERXSTATUSL6,
    PIPERXSTATUSL7,
    PIPERXVALIDL0,
    PIPERXVALIDL1,
    PIPERXVALIDL2,
    PIPERXVALIDL3,
    PIPERXVALIDL4,
    PIPERXVALIDL5,
    PIPERXVALIDL6,
    PIPERXVALIDL7

);

parameter AERCAPABILITYECRCCHECKCAPABLE = "FALSE";
parameter AERCAPABILITYECRCGENCAPABLE = "FALSE";
parameter BAR0EXIST = "TRUE";
parameter BAR0PREFETCHABLE = "TRUE";
parameter BAR1EXIST = "FALSE";
parameter BAR1PREFETCHABLE = "FALSE";
parameter BAR2EXIST = "FALSE";
parameter BAR2PREFETCHABLE = "FALSE";
parameter BAR3EXIST = "FALSE";
parameter BAR3PREFETCHABLE = "FALSE";
parameter BAR4EXIST = "FALSE";
parameter BAR4PREFETCHABLE = "FALSE";
parameter BAR5EXIST = "FALSE";
parameter BAR5PREFETCHABLE = "FALSE";
parameter CLKDIVIDED = "FALSE";
parameter DUALCOREENABLE = "FALSE";
parameter DUALCORESLAVE = "FALSE";
parameter INFINITECOMPLETIONS = "TRUE";
parameter ISSWITCH = "FALSE";
parameter LINKSTATUSSLOTCLOCKCONFIG = "FALSE";
parameter LLKBYPASS = "FALSE";
parameter PBCAPABILITYSYSTEMALLOCATED = "FALSE";
parameter PCIECAPABILITYSLOTIMPL = "FALSE";
parameter PMCAPABILITYD1SUPPORT = "FALSE";
parameter PMCAPABILITYD2SUPPORT = "FALSE";
parameter PMCAPABILITYDSI = "TRUE";
parameter RAMSHARETXRX = "FALSE";
parameter RESETMODE = "FALSE";
parameter RETRYREADADDRPIPE = "FALSE";
parameter RETRYREADDATAPIPE = "FALSE";
parameter RETRYWRITEPIPE = "FALSE";
parameter RXREADADDRPIPE = "FALSE";
parameter RXREADDATAPIPE = "FALSE";
parameter RXWRITEPIPE = "FALSE";
parameter SELECTASMODE = "FALSE";
parameter SELECTDLLIF = "FALSE";
parameter SLOTCAPABILITYATTBUTTONPRESENT = "FALSE";
parameter SLOTCAPABILITYATTINDICATORPRESENT = "FALSE";
parameter SLOTCAPABILITYHOTPLUGCAPABLE = "FALSE";
parameter SLOTCAPABILITYHOTPLUGSURPRISE = "FALSE";
parameter SLOTCAPABILITYMSLSENSORPRESENT = "FALSE";
parameter SLOTCAPABILITYPOWERCONTROLLERPRESENT = "FALSE";
parameter SLOTCAPABILITYPOWERINDICATORPRESENT = "FALSE";
parameter SLOTIMPLEMENTED = "FALSE";
parameter TXREADADDRPIPE = "FALSE";
parameter TXREADDATAPIPE = "FALSE";
parameter TXWRITEPIPE = "FALSE";
parameter UPSTREAMFACING = "TRUE";
parameter XLINKSUPPORTED = "FALSE";
parameter [10:0] VC0TOTALCREDITSCD = 11'h0;
parameter [10:0] VC0TOTALCREDITSPD = 11'h34;
parameter [10:0] VC1TOTALCREDITSCD = 11'h0;
parameter [10:0] VC1TOTALCREDITSPD = 11'h0;
parameter [11:0] AERBASEPTR = 12'h110;
parameter [11:0] AERCAPABILITYNEXTPTR = 12'h138;
parameter [11:0] DSNBASEPTR = 12'h148;
parameter [11:0] DSNCAPABILITYNEXTPTR = 12'h154;
parameter [11:0] EXTCFGXPCAPPTR = 12'h0;
parameter [11:0] MSIBASEPTR = 12'h48;
parameter [11:0] PBBASEPTR = 12'h138;
parameter [11:0] PBCAPABILITYNEXTPTR = 12'h148;
parameter [11:0] PMBASEPTR = 12'h40;
parameter [11:0] RETRYRAMSIZE = 12'h9;
parameter [11:0] VCBASEPTR = 12'h154;
parameter [11:0] VCCAPABILITYNEXTPTR = 12'h0;
parameter [12:0] SLOTCAPABILITYPHYSICALSLOTNUM = 13'h0;
parameter [12:0] VC0RXFIFOBASEC = 13'h98;
parameter [12:0] VC0RXFIFOBASENP = 13'h80;
parameter [12:0] VC0RXFIFOBASEP = 13'h0;
parameter [12:0] VC0RXFIFOLIMITC = 13'h117;
parameter [12:0] VC0RXFIFOLIMITNP = 13'h97;
parameter [12:0] VC0RXFIFOLIMITP = 13'h7f;
parameter [12:0] VC0TXFIFOBASEC = 13'h98;
parameter [12:0] VC0TXFIFOBASENP = 13'h80;
parameter [12:0] VC0TXFIFOBASEP = 13'h0;
parameter [12:0] VC0TXFIFOLIMITC = 13'h117;
parameter [12:0] VC0TXFIFOLIMITNP = 13'h97;
parameter [12:0] VC0TXFIFOLIMITP = 13'h7f;
parameter [12:0] VC1RXFIFOBASEC = 13'h118;
parameter [12:0] VC1RXFIFOBASENP = 13'h118;
parameter [12:0] VC1RXFIFOBASEP = 13'h118;
parameter [12:0] VC1RXFIFOLIMITC = 13'h118;
parameter [12:0] VC1RXFIFOLIMITNP = 13'h118;
parameter [12:0] VC1RXFIFOLIMITP = 13'h118;
parameter [12:0] VC1TXFIFOBASEC = 13'h118;
parameter [12:0] VC1TXFIFOBASENP = 13'h118;
parameter [12:0] VC1TXFIFOBASEP = 13'h118;
parameter [12:0] VC1TXFIFOLIMITC = 13'h118;
parameter [12:0] VC1TXFIFOLIMITNP = 13'h118;
parameter [12:0] VC1TXFIFOLIMITP = 13'h118;
parameter [15:0] DEVICEID = 16'h5050;
parameter [15:0] SUBSYSTEMID = 16'h5050;
parameter [15:0] SUBSYSTEMVENDORID = 16'h10EE;
parameter [15:0] VENDORID = 16'h10EE;
parameter [1:0] LINKCAPABILITYASPMSUPPORT = 2'h1;
parameter [1:0] PBCAPABILITYDW0DATASCALE = 2'h0;
parameter [1:0] PBCAPABILITYDW0PMSTATE = 2'h0;
parameter [1:0] PBCAPABILITYDW1DATASCALE = 2'h0;
parameter [1:0] PBCAPABILITYDW1PMSTATE = 2'h0;
parameter [1:0] PBCAPABILITYDW2DATASCALE = 2'h0;
parameter [1:0] PBCAPABILITYDW2PMSTATE = 2'h0;
parameter [1:0] PBCAPABILITYDW3DATASCALE = 2'h0;
parameter [1:0] PBCAPABILITYDW3PMSTATE = 2'h0;
parameter [1:0] PMSTATUSCONTROLDATASCALE = 2'h0;
parameter [1:0] SLOTCAPABILITYSLOTPOWERLIMITSCALE = 2'h0;
parameter [23:0] CLASSCODE = 24'h058000;
parameter [2:0] CONFIGROUTING = 3'h1;
parameter [2:0] DEVICECAPABILITYENDPOINTL0SLATENCY = 3'h0;
parameter [2:0] DEVICECAPABILITYENDPOINTL1LATENCY = 3'h0;
parameter [2:0] MSICAPABILITYMULTIMSGCAP = 3'h0;
parameter [2:0] PBCAPABILITYDW0PMSUBSTATE = 3'h0;
parameter [2:0] PBCAPABILITYDW0POWERRAIL = 3'h0;
parameter [2:0] PBCAPABILITYDW0TYPE = 3'h0;
parameter [2:0] PBCAPABILITYDW1PMSUBSTATE = 3'h0;
parameter [2:0] PBCAPABILITYDW1POWERRAIL = 3'h0;
parameter [2:0] PBCAPABILITYDW1TYPE = 3'h0;
parameter [2:0] PBCAPABILITYDW2PMSUBSTATE = 3'h0;
parameter [2:0] PBCAPABILITYDW2POWERRAIL = 3'h0;
parameter [2:0] PBCAPABILITYDW2TYPE = 3'h0;
parameter [2:0] PBCAPABILITYDW3PMSUBSTATE = 3'h0;
parameter [2:0] PBCAPABILITYDW3POWERRAIL = 3'h0;
parameter [2:0] PBCAPABILITYDW3TYPE = 3'h0;
parameter [2:0] PMCAPABILITYAUXCURRENT = 3'h0;
parameter [2:0] PORTVCCAPABILITYEXTENDEDVCCOUNT = 3'h0;
parameter [31:0] CARDBUSCISPOINTER = 32'h0;
parameter [3:0] XPDEVICEPORTTYPE = 4'h0;
parameter [4:0] PCIECAPABILITYINTMSGNUM = 5'h0;
parameter [4:0] PMCAPABILITYPMESUPPORT = 5'h0;
parameter [5:0] BAR0MASKWIDTH = 6'h14;
parameter [5:0] BAR1MASKWIDTH = 6'h0;
parameter [5:0] BAR2MASKWIDTH = 6'h0;
parameter [5:0] BAR3MASKWIDTH = 6'h0;
parameter [5:0] BAR4MASKWIDTH = 6'h0;
parameter [5:0] BAR5MASKWIDTH = 6'h0;
parameter [5:0] LINKCAPABILITYMAXLINKWIDTH = 6'h01;
parameter [63:0] DEVICESERIALNUMBER = 64'hE000000001000A35;
parameter [6:0] VC0TOTALCREDITSCH = 7'h0;
parameter [6:0] VC0TOTALCREDITSNPH = 7'h08;
parameter [6:0] VC0TOTALCREDITSPH = 7'h08;
parameter [6:0] VC1TOTALCREDITSCH = 7'h0;
parameter [6:0] VC1TOTALCREDITSNPH = 7'h0;
parameter [6:0] VC1TOTALCREDITSPH = 7'h0;
parameter [7:0] ACTIVELANESIN = 8'h1;
parameter [7:0] CAPABILITIESPOINTER = 8'h40;
parameter [7:0] EXTCFGCAPPTR = 8'h0;
parameter [7:0] HEADERTYPE = 8'h0;
parameter [7:0] INTERRUPTPIN = 8'h0;
parameter [7:0] MSICAPABILITYNEXTPTR = 8'h60;
parameter [7:0] PBCAPABILITYDW0BASEPOWER = 8'h0;
parameter [7:0] PBCAPABILITYDW1BASEPOWER = 8'h0;
parameter [7:0] PBCAPABILITYDW2BASEPOWER = 8'h0;
parameter [7:0] PBCAPABILITYDW3BASEPOWER = 8'h0;
parameter [7:0] PCIECAPABILITYNEXTPTR = 8'h0;
parameter [7:0] PMCAPABILITYNEXTPTR = 8'h60;
parameter [7:0] PMDATA0 = 8'h0;
parameter [7:0] PMDATA1 = 8'h0;
parameter [7:0] PMDATA2 = 8'h0;
parameter [7:0] PMDATA3 = 8'h0;
parameter [7:0] PMDATA4 = 8'h0;
parameter [7:0] PMDATA5 = 8'h0;
parameter [7:0] PMDATA6 = 8'h0;
parameter [7:0] PMDATA7 = 8'h0;
parameter [7:0] PMDATA8 = 8'h0;
parameter [7:0] PORTVCCAPABILITYVCARBCAP = 8'h0;
parameter [7:0] PORTVCCAPABILITYVCARBTABLEOFFSET = 8'h0;
parameter [7:0] REVISIONID = 8'h0;
parameter [7:0] SLOTCAPABILITYSLOTPOWERLIMITVALUE = 8'h0;
parameter [7:0] XPBASEPTR = 8'h60;
parameter BAR0ADDRWIDTH = 0;
parameter BAR0IOMEMN = 0;
parameter BAR1ADDRWIDTH = 0;
parameter BAR1IOMEMN = 0;
parameter BAR2ADDRWIDTH = 0;
parameter BAR2IOMEMN = 0;
parameter BAR3ADDRWIDTH = 0;
parameter BAR3IOMEMN = 0;
parameter BAR4ADDRWIDTH = 0;
parameter BAR4IOMEMN = 0;
parameter BAR5IOMEMN = 0;
parameter DUALROLECFGCNTRLROOTEPN = 0;
parameter L0SEXITLATENCY = 7;
parameter L0SEXITLATENCYCOMCLK = 7;
parameter L1EXITLATENCY = 7;
parameter L1EXITLATENCYCOMCLK = 7;
parameter LOWPRIORITYVCCOUNT = 0;
parameter PCIEREVISION = 1;
parameter PMDATASCALE0 = 0;
parameter PMDATASCALE1 = 0;
parameter PMDATASCALE2 = 0;
parameter PMDATASCALE3 = 0;
parameter PMDATASCALE4 = 0;
parameter PMDATASCALE5 = 0;
parameter PMDATASCALE6 = 0;
parameter PMDATASCALE7 = 0;
parameter PMDATASCALE8 = 0;
parameter RETRYRAMREADLATENCY = 3;
parameter RETRYRAMWIDTH = 0;
parameter RETRYRAMWRITELATENCY = 1;
parameter TLRAMREADLATENCY = 3;
parameter TLRAMWIDTH = 0;
parameter TLRAMWRITELATENCY = 1;
parameter TXTSNFTS = 255;
parameter TXTSNFTSCOMCLK = 255;
parameter XPMAXPAYLOAD = 0;
parameter XPRCBCONTROL = 0;


output BUSMASTERENABLE;
output CRMDOHOTRESETN;
output CRMPWRSOFTRESETN;
output CRMRXHOTRESETN;
output DLLTXPMDLLPOUTSTANDING;
output INTERRUPTDISABLE;
output IOSPACEENABLE;
output L0ASAUTONOMOUSINITCOMPLETED;
output L0CFGLOOPBACKACK;
output L0CORRERRMSGRCVD;
output L0DLLASTXSTATE;
output L0DLLRXACKOUTSTANDING;
output L0DLLTXNONFCOUTSTANDING;
output L0DLLTXOUTSTANDING;
output L0FATALERRMSGRCVD;
output L0FIRSTCFGWRITEOCCURRED;
output L0FWDCORRERROUT;
output L0FWDFATALERROUT;
output L0FWDNONFATALERROUT;
output L0MACENTEREDL0;
output L0MACLINKTRAINING;
output L0MACLINKUP;
output L0MACNEWSTATEACK;
output L0MACRXL0SSTATE;
output L0MACUPSTREAMDOWNSTREAM;
output L0MSIENABLE0;
output L0NONFATALERRMSGRCVD;
output L0PMEACK;
output L0PMEEN;
output L0PMEREQOUT;
output L0POWERCONTROLLERCONTROL;
output L0PWRINHIBITTRANSFERS;
output L0PWRL1STATE;
output L0PWRL23READYDEVICE;
output L0PWRL23READYSTATE;
output L0PWRTURNOFFREQ;
output L0PWRTXL0SSTATE;
output L0RECEIVEDASSERTINTALEGACYINT;
output L0RECEIVEDASSERTINTBLEGACYINT;
output L0RECEIVEDASSERTINTCLEGACYINT;
output L0RECEIVEDASSERTINTDLEGACYINT;
output L0RECEIVEDDEASSERTINTALEGACYINT;
output L0RECEIVEDDEASSERTINTBLEGACYINT;
output L0RECEIVEDDEASSERTINTCLEGACYINT;
output L0RECEIVEDDEASSERTINTDLEGACYINT;
output L0RXBEACON;
output L0RXDLLPM;
output L0RXDLLSBFCUPDATE;
output L0RXDLLTLPECRCOK;
output L0STATSCFGOTHERRECEIVED;
output L0STATSCFGOTHERTRANSMITTED;
output L0STATSCFGRECEIVED;
output L0STATSCFGTRANSMITTED;
output L0STATSDLLPRECEIVED;
output L0STATSDLLPTRANSMITTED;
output L0STATSOSRECEIVED;
output L0STATSOSTRANSMITTED;
output L0STATSTLPRECEIVED;
output L0STATSTLPTRANSMITTED;
output L0TOGGLEELECTROMECHANICALINTERLOCK;
output L0TXDLLPMUPDATED;
output L0TXDLLSBFCUPDATED;
output L0UNLOCKRECEIVED;
output LLKRX4DWHEADERN;
output LLKRXCHCONFIGAVAILABLEN;
output LLKRXCHCONFIGPARTIALN;
output LLKRXECRCBADN;
output LLKRXEOFN;
output LLKRXEOPN;
output LLKRXSOFN;
output LLKRXSOPN;
output LLKRXSRCDSCN;
output LLKRXSRCLASTREQN;
output LLKRXSRCRDYN;
output LLKTXCONFIGREADYN;
output LLKTXDSTRDYN;
output MEMSPACEENABLE;
output MIMDLLBREN;
output MIMDLLBWEN;
output MIMRXBREN;
output MIMRXBWEN;
output MIMTXBREN;
output MIMTXBWEN;
output PARITYERRORRESPONSE;
output PIPEDESKEWLANESL0;
output PIPEDESKEWLANESL1;
output PIPEDESKEWLANESL2;
output PIPEDESKEWLANESL3;
output PIPEDESKEWLANESL4;
output PIPEDESKEWLANESL5;
output PIPEDESKEWLANESL6;
output PIPEDESKEWLANESL7;
output PIPERESETL0;
output PIPERESETL1;
output PIPERESETL2;
output PIPERESETL3;
output PIPERESETL4;
output PIPERESETL5;
output PIPERESETL6;
output PIPERESETL7;
output PIPERXPOLARITYL0;
output PIPERXPOLARITYL1;
output PIPERXPOLARITYL2;
output PIPERXPOLARITYL3;
output PIPERXPOLARITYL4;
output PIPERXPOLARITYL5;
output PIPERXPOLARITYL6;
output PIPERXPOLARITYL7;
output PIPETXCOMPLIANCEL0;
output PIPETXCOMPLIANCEL1;
output PIPETXCOMPLIANCEL2;
output PIPETXCOMPLIANCEL3;
output PIPETXCOMPLIANCEL4;
output PIPETXCOMPLIANCEL5;
output PIPETXCOMPLIANCEL6;
output PIPETXCOMPLIANCEL7;
output PIPETXDATAKL0;
output PIPETXDATAKL1;
output PIPETXDATAKL2;
output PIPETXDATAKL3;
output PIPETXDATAKL4;
output PIPETXDATAKL5;
output PIPETXDATAKL6;
output PIPETXDATAKL7;
output PIPETXDETECTRXLOOPBACKL0;
output PIPETXDETECTRXLOOPBACKL1;
output PIPETXDETECTRXLOOPBACKL2;
output PIPETXDETECTRXLOOPBACKL3;
output PIPETXDETECTRXLOOPBACKL4;
output PIPETXDETECTRXLOOPBACKL5;
output PIPETXDETECTRXLOOPBACKL6;
output PIPETXDETECTRXLOOPBACKL7;
output PIPETXELECIDLEL0;
output PIPETXELECIDLEL1;
output PIPETXELECIDLEL2;
output PIPETXELECIDLEL3;
output PIPETXELECIDLEL4;
output PIPETXELECIDLEL5;
output PIPETXELECIDLEL6;
output PIPETXELECIDLEL7;
output SERRENABLE;
output URREPORTINGENABLE;
output [11:0] MGMTSTATSCREDIT;
output [11:0] MIMDLLBRADD;
output [11:0] MIMDLLBWADD;
output [12:0] L0COMPLETERID;
output [12:0] MIMRXBRADD;
output [12:0] MIMRXBWADD;
output [12:0] MIMTXBRADD;
output [12:0] MIMTXBWADD;
output [15:0] L0ERRMSGREQID;
output [15:0] LLKRXPREFERREDTYPE;
output [16:0] MGMTPSO;
output [18:0] L0RXDLLSBFCDATA;
output [19:0] L0RXDLLFCNPOSTBYPCRED;
output [1:0] L0ATTENTIONINDICATORCONTROL;
output [1:0] L0DLLASRXSTATE;
output [1:0] L0POWERINDICATORCONTROL;
output [1:0] L0PWRSTATE0;
output [1:0] L0RXDLLTLPEND;
output [1:0] L0RXMACLINKERROR;
output [1:0] LLKRXVALIDN;
output [1:0] PIPEPOWERDOWNL0;
output [1:0] PIPEPOWERDOWNL1;
output [1:0] PIPEPOWERDOWNL2;
output [1:0] PIPEPOWERDOWNL3;
output [1:0] PIPEPOWERDOWNL4;
output [1:0] PIPEPOWERDOWNL5;
output [1:0] PIPEPOWERDOWNL6;
output [1:0] PIPEPOWERDOWNL7;
output [23:0] L0RXDLLFCCMPLMCCRED;
output [23:0] L0RXDLLFCPOSTORDCRED;
output [2:0] L0MCFOUND;
output [2:0] L0MULTIMSGEN0;
output [2:0] L0RXDLLPMTYPE;
output [2:0] L0TRANSFORMEDVC;
output [2:0] MAXPAYLOADSIZE;
output [2:0] MAXREADREQUESTSIZE;
output [31:0] MGMTRDATA;
output [3:0] L0LTSSMSTATE;
output [3:0] L0MACNEGOTIATEDLINKWIDTH;
output [3:0] L0UCBYPFOUND;
output [3:0] L0UCORDFOUND;
output [63:0] LLKRXDATA;
output [63:0] MIMDLLBWDATA;
output [63:0] MIMRXBWDATA;
output [63:0] MIMTXBWDATA;
output [6:0] L0DLLERRORVECTOR;
output [7:0] L0DLLVCSTATUS;
output [7:0] L0DLUPDOWN;
output [7:0] L0RXDLLFCCMPLMCUPDATE;
output [7:0] L0RXDLLFCNPOSTBYPUPDATE;
output [7:0] L0RXDLLFCPOSTORDUPDATE;
output [7:0] L0TXDLLFCCMPLMCUPDATED;
output [7:0] L0TXDLLFCNPOSTBYPUPDATED;
output [7:0] L0TXDLLFCPOSTORDUPDATED;
output [7:0] LLKRXCHCOMPLETIONAVAILABLEN;
output [7:0] LLKRXCHCOMPLETIONPARTIALN;
output [7:0] LLKRXCHNONPOSTEDAVAILABLEN;
output [7:0] LLKRXCHNONPOSTEDPARTIALN;
output [7:0] LLKRXCHPOSTEDAVAILABLEN;
output [7:0] LLKRXCHPOSTEDPARTIALN;
output [7:0] LLKTCSTATUS;
output [7:0] LLKTXCHCOMPLETIONREADYN;
output [7:0] LLKTXCHNONPOSTEDREADYN;
output [7:0] LLKTXCHPOSTEDREADYN;
output [7:0] PIPETXDATAL0;
output [7:0] PIPETXDATAL1;
output [7:0] PIPETXDATAL2;
output [7:0] PIPETXDATAL3;
output [7:0] PIPETXDATAL4;
output [7:0] PIPETXDATAL5;
output [7:0] PIPETXDATAL6;
output [7:0] PIPETXDATAL7;
output [9:0] LLKTXCHANSPACE;

input AUXPOWER;
input COMPLIANCEAVOID;
input CRMCFGBRIDGEHOTRESET;
input CRMCORECLK;
input CRMCORECLKDLO;
input CRMCORECLKRXO;
input CRMCORECLKTXO;
input CRMLINKRSTN;
input CRMMACRSTN;
input CRMMGMTRSTN;
input CRMNVRSTN;
input CRMTXHOTRESETN;
input CRMURSTN;
input CRMUSERCFGRSTN;
input CRMUSERCLK;
input CRMUSERCLKRXO;
input CRMUSERCLKTXO;
input CROSSLINKSEED;
input L0ALLDOWNPORTSINL1;
input L0ALLDOWNRXPORTSINL0S;
input L0ASE;
input L0ATTENTIONBUTTONPRESSED;
input L0CFGASSPANTREEOWNEDSTATE;
input L0CFGDISABLESCRAMBLE;
input L0CFGEXTENDEDSYNC;
input L0CFGL0SENTRYENABLE;
input L0CFGL0SENTRYSUP;
input L0CFGLINKDISABLE;
input L0CFGLOOPBACKMASTER;
input L0DLLHOLDLINKUP;
input L0ELECTROMECHANICALINTERLOCKENGAGED;
input L0FWDASSERTINTALEGACYINT;
input L0FWDASSERTINTBLEGACYINT;
input L0FWDASSERTINTCLEGACYINT;
input L0FWDASSERTINTDLEGACYINT;
input L0FWDCORRERRIN;
input L0FWDDEASSERTINTALEGACYINT;
input L0FWDDEASSERTINTBLEGACYINT;
input L0FWDDEASSERTINTCLEGACYINT;
input L0FWDDEASSERTINTDLEGACYINT;
input L0FWDFATALERRIN;
input L0FWDNONFATALERRIN;
input L0LEGACYINTFUNCT0;
input L0MRLSENSORCLOSEDN;
input L0PMEREQIN;
input L0POWERFAULTDETECTED;
input L0PRESENCEDETECTSLOTEMPTYN;
input L0PWRNEWSTATEREQ;
input L0ROOTTURNOFFREQ;
input L0SENDUNLOCKMESSAGE;
input L0SETCOMPLETERABORTERROR;
input L0SETCOMPLETIONTIMEOUTCORRERROR;
input L0SETCOMPLETIONTIMEOUTUNCORRERROR;
input L0SETDETECTEDCORRERROR;
input L0SETDETECTEDFATALERROR;
input L0SETDETECTEDNONFATALERROR;
input L0SETLINKDETECTEDPARITYERROR;
input L0SETLINKMASTERDATAPARITY;
input L0SETLINKRECEIVEDMASTERABORT;
input L0SETLINKRECEIVEDTARGETABORT;
input L0SETLINKSIGNALLEDTARGETABORT;
input L0SETLINKSYSTEMERROR;
input L0SETUNEXPECTEDCOMPLETIONCORRERROR;
input L0SETUNEXPECTEDCOMPLETIONUNCORRERROR;
input L0SETUNSUPPORTEDREQUESTNONPOSTEDERROR;
input L0SETUNSUPPORTEDREQUESTOTHERERROR;
input L0SETUSERDETECTEDPARITYERROR;
input L0SETUSERMASTERDATAPARITY;
input L0SETUSERRECEIVEDMASTERABORT;
input L0SETUSERRECEIVEDTARGETABORT;
input L0SETUSERSIGNALLEDTARGETABORT;
input L0SETUSERSYSTEMERROR;
input L0TLASFCCREDSTARVATION;
input L0TLLINKRETRAIN;
input L0TRANSACTIONSPENDING;
input L0TXBEACON;
input L0TXCFGPM;
input L0TXTLSBFCUPDATE;
input L0TXTLTLPEDB;
input L0TXTLTLPREQ;
input L0TXTLTLPREQEND;
input L0TXTLTLPWIDTH;
input L0UPSTREAMRXPORTINL0S;
input L0VC0PREVIEWEXPAND;
input L0WAKEN;
input LLKRXDSTCONTREQN;
input LLKRXDSTREQN;
input LLKTX4DWHEADERN;
input LLKTXCOMPLETEN;
input LLKTXCREATEECRCN;
input LLKTXEOFN;
input LLKTXEOPN;
input LLKTXSOFN;
input LLKTXSOPN;
input LLKTXSRCDSCN;
input LLKTXSRCRDYN;
input MAINPOWER;
input MGMTRDEN;
input MGMTWREN;
input PIPEPHYSTATUSL0;
input PIPEPHYSTATUSL1;
input PIPEPHYSTATUSL2;
input PIPEPHYSTATUSL3;
input PIPEPHYSTATUSL4;
input PIPEPHYSTATUSL5;
input PIPEPHYSTATUSL6;
input PIPEPHYSTATUSL7;
input PIPERXCHANISALIGNEDL0;
input PIPERXCHANISALIGNEDL1;
input PIPERXCHANISALIGNEDL2;
input PIPERXCHANISALIGNEDL3;
input PIPERXCHANISALIGNEDL4;
input PIPERXCHANISALIGNEDL5;
input PIPERXCHANISALIGNEDL6;
input PIPERXCHANISALIGNEDL7;
input PIPERXDATAKL0;
input PIPERXDATAKL1;
input PIPERXDATAKL2;
input PIPERXDATAKL3;
input PIPERXDATAKL4;
input PIPERXDATAKL5;
input PIPERXDATAKL6;
input PIPERXDATAKL7;
input PIPERXELECIDLEL0;
input PIPERXELECIDLEL1;
input PIPERXELECIDLEL2;
input PIPERXELECIDLEL3;
input PIPERXELECIDLEL4;
input PIPERXELECIDLEL5;
input PIPERXELECIDLEL6;
input PIPERXELECIDLEL7;
input PIPERXVALIDL0;
input PIPERXVALIDL1;
input PIPERXVALIDL2;
input PIPERXVALIDL3;
input PIPERXVALIDL4;
input PIPERXVALIDL5;
input PIPERXVALIDL6;
input PIPERXVALIDL7;
input [10:0] MGMTADDR;
input [11:0] L0ACKNAKTIMERADJUSTMENT;
input [11:0] L0REPLAYTIMERADJUSTMENT;
input [127:0] L0PACKETHEADERFROMUSER;
input [159:0] L0TXTLFCCMPLMCCRED;
input [159:0] L0TXTLFCPOSTORDCRED;
input [15:0] L0TXTLFCCMPLMCUPDATE;
input [15:0] L0TXTLFCNPOSTBYPUPDATE;
input [15:0] L0TXTLFCPOSTORDUPDATE;
input [18:0] L0TXTLSBFCDATA;
input [191:0] L0TXTLFCNPOSTBYPCRED;
input [1:0] L0PWRNEXTLINKSTATE;
input [1:0] L0TXTLTLPENABLE;
input [1:0] L0TXTLTLPEND;
input [1:0] LLKRXCHFIFO;
input [1:0] LLKTXCHFIFO;
input [1:0] LLKTXENABLEN;
input [23:0] L0CFGVCID;
input [2:0] L0ASTURNPOOLBITSCONSUMED;
input [2:0] L0CFGL0SEXITLAT;
input [2:0] L0CFGNEGOTIATEDMAXP;
input [2:0] L0TXCFGPMTYPE;
input [2:0] LLKRXCHTC;
input [2:0] LLKTXCHTC;
input [2:0] PIPERXSTATUSL0;
input [2:0] PIPERXSTATUSL1;
input [2:0] PIPERXSTATUSL2;
input [2:0] PIPERXSTATUSL3;
input [2:0] PIPERXSTATUSL4;
input [2:0] PIPERXSTATUSL5;
input [2:0] PIPERXSTATUSL6;
input [2:0] PIPERXSTATUSL7;
input [31:0] MGMTWDATA;
input [3:0] L0CFGASSTATECHANGECMD;
input [3:0] L0MSIREQUEST0;
input [3:0] L0TXTLTLPLATENCY;
input [3:0] MGMTBWREN;
input [5:0] CFGNEGOTIATEDLINKWIDTH;
input [63:0] L0TXTLTLPDATA;
input [63:0] LLKTXDATA;
input [63:0] MIMDLLBRDATA;
input [63:0] MIMRXBRDATA;
input [63:0] MIMTXBRDATA;
input [6:0] MGMTSTATSCREDITSEL;
input [7:0] L0ASPORTCOUNT;
input [7:0] L0CFGVCENABLE;
input [7:0] L0PORTNUMBER;
input [7:0] L0RXTLTLPNONINITIALIZEDVC;
input [7:0] PIPERXDATAL0;
input [7:0] PIPERXDATAL1;
input [7:0] PIPERXDATAL2;
input [7:0] PIPERXDATAL3;
input [7:0] PIPERXDATAL4;
input [7:0] PIPERXDATAL5;
input [7:0] PIPERXDATAL6;
input [7:0] PIPERXDATAL7;

endmodule
