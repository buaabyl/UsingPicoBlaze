///////////////////////////////////////////////////////
//  Copyright (c) 2008 Xilinx Inc.
//  All Right Reserved.
///////////////////////////////////////////////////////
//
//   ____   ___
//  /   /\/   / 
// /___/  \  /     Vendor      : Xilinx 
// \  \    \/      Version     : 12.i 
//  \  \           Description : 
//  /  /                      
// /__/   /\       Filename    : X_POST_CRC_INTERNAL.v
// \  \  /  \ 
//  \__\/\__ \                    
//                                 
//  Revision:        1.0
///////////////////////////////////////////////////////

`timescale 1 ps / 1 ps 

module X_POST_CRC_INTERNAL (
  CRCERROR
);

  output CRCERROR;
 
endmodule
