//    Xilinx Proprietary Primitive Cell X_IPAD for Verilog
//
// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/xec_libs/data/simprims/X_IPAD.v,v 1.2 2008/10/02 19:01:54 vandanad Exp $
//

`celldefine
`timescale 1 ps/1 ps

module X_IPAD (PAD);

  input PAD;
  parameter LOC = "UNPLACED";
endmodule
