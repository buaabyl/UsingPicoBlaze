//    Xilinx Proprietary Primitive Cell X_SUH for Verilog
//
// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/xec_libs/data/simprims/X_SUH.v,v 1.2 2008/10/02 19:01:56 vandanad Exp $
//

`celldefine
`timescale 1 ps/1 ps

module X_SUH (I, CE, CLK);

  input I, CLK, CE;
  parameter LOC = "UNPLACED";
endmodule
