// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/xec_libs/data/simprims/X_EMAC.v,v 1.2 2008/10/02 19:01:53 vandanad Exp $

`timescale 1 ps / 1 ps 

module X_EMAC (
    DCRHOSTDONEIR,
    EMAC0CLIENTANINTERRUPT,
    EMAC0CLIENTRXBADFRAME,
    EMAC0CLIENTRXCLIENTCLKOUT,
    EMAC0CLIENTRXD,
    EMAC0CLIENTRXDVLD,
    EMAC0CLIENTRXDVLDMSW,
    EMAC0CLIENTRXDVREG6,
    EMAC0CLIENTRXFRAMEDROP,
    EMAC0CLIENTRXGOODFRAME,
    EMAC0CLIENTRXSTATS,
    EMAC0CLIENTRXSTATSBYTEVLD,
    EMAC0CLIENTRXSTATSVLD,
    EMAC0CLIENTTXACK,
    EMAC0CLIENTTXCLIENTCLKOUT,
    EMAC0CLIENTTXCOLLISION,
    EMAC0CLIENTTXGMIIMIICLKOUT,
    EMAC0CLIENTTXRETRANSMIT,
    EMAC0CLIENTTXSTATS,
    EMAC0CLIENTTXSTATSBYTEVLD,
    EMAC0CLIENTTXSTATSVLD,
    EMAC0PHYENCOMMAALIGN,
    EMAC0PHYLOOPBACKMSB,
    EMAC0PHYMCLKOUT,
    EMAC0PHYMDOUT,
    EMAC0PHYMDTRI,
    EMAC0PHYMGTRXRESET,
    EMAC0PHYMGTTXRESET,
    EMAC0PHYPOWERDOWN,
    EMAC0PHYSYNCACQSTATUS,
    EMAC0PHYTXCHARDISPMODE,
    EMAC0PHYTXCHARDISPVAL,
    EMAC0PHYTXCHARISK,
    EMAC0PHYTXCLK,
    EMAC0PHYTXD,
    EMAC0PHYTXEN,
    EMAC0PHYTXER,
    EMAC1CLIENTANINTERRUPT,
    EMAC1CLIENTRXBADFRAME,
    EMAC1CLIENTRXCLIENTCLKOUT,
    EMAC1CLIENTRXD,
    EMAC1CLIENTRXDVLD,
    EMAC1CLIENTRXDVLDMSW,
    EMAC1CLIENTRXDVREG6,
    EMAC1CLIENTRXFRAMEDROP,
    EMAC1CLIENTRXGOODFRAME,
    EMAC1CLIENTRXSTATS,
    EMAC1CLIENTRXSTATSBYTEVLD,
    EMAC1CLIENTRXSTATSVLD,
    EMAC1CLIENTTXACK,
    EMAC1CLIENTTXCLIENTCLKOUT,
    EMAC1CLIENTTXCOLLISION,
    EMAC1CLIENTTXGMIIMIICLKOUT,
    EMAC1CLIENTTXRETRANSMIT,
    EMAC1CLIENTTXSTATS,
    EMAC1CLIENTTXSTATSBYTEVLD,
    EMAC1CLIENTTXSTATSVLD,
    EMAC1PHYENCOMMAALIGN,
    EMAC1PHYLOOPBACKMSB,
    EMAC1PHYMCLKOUT,
    EMAC1PHYMDOUT,
    EMAC1PHYMDTRI,
    EMAC1PHYMGTRXRESET,
    EMAC1PHYMGTTXRESET,
    EMAC1PHYPOWERDOWN,
    EMAC1PHYSYNCACQSTATUS,
    EMAC1PHYTXCHARDISPMODE,
    EMAC1PHYTXCHARDISPVAL,
    EMAC1PHYTXCHARISK,
    EMAC1PHYTXCLK,
    EMAC1PHYTXD,
    EMAC1PHYTXEN,
    EMAC1PHYTXER,
    EMACDCRACK,
    EMACDCRDBUS,
    HOSTMIIMRDY,
    HOSTRDDATA,
    CLIENTEMAC0DCMLOCKED,
    CLIENTEMAC0PAUSEREQ,
    CLIENTEMAC0PAUSEVAL,
    CLIENTEMAC0RXCLIENTCLKIN,
    CLIENTEMAC0TXCLIENTCLKIN,
    CLIENTEMAC0TXD,
    CLIENTEMAC0TXDVLD,
    CLIENTEMAC0TXDVLDMSW,
    CLIENTEMAC0TXFIRSTBYTE,
    CLIENTEMAC0TXGMIIMIICLKIN,
    CLIENTEMAC0TXIFGDELAY,
    CLIENTEMAC0TXUNDERRUN,
    CLIENTEMAC1DCMLOCKED,
    CLIENTEMAC1PAUSEREQ,
    CLIENTEMAC1PAUSEVAL,
    CLIENTEMAC1RXCLIENTCLKIN,
    CLIENTEMAC1TXCLIENTCLKIN,
    CLIENTEMAC1TXD,
    CLIENTEMAC1TXDVLD,
    CLIENTEMAC1TXDVLDMSW,
    CLIENTEMAC1TXFIRSTBYTE,
    CLIENTEMAC1TXGMIIMIICLKIN,
    CLIENTEMAC1TXIFGDELAY,
    CLIENTEMAC1TXUNDERRUN,
    DCREMACABUS,
    DCREMACCLK,
    DCREMACDBUS,
    DCREMACENABLE,
    DCREMACREAD,
    DCREMACWRITE,
    HOSTADDR,
    HOSTCLK,
    HOSTEMAC1SEL,
    HOSTMIIMSEL,
    HOSTOPCODE,
    HOSTREQ,
    HOSTWRDATA,
    PHYEMAC0COL,
    PHYEMAC0CRS,
    PHYEMAC0GTXCLK,
    PHYEMAC0MCLKIN,
    PHYEMAC0MDIN,
    PHYEMAC0MIITXCLK,
    PHYEMAC0PHYAD,
    PHYEMAC0RXBUFERR,
    PHYEMAC0RXBUFSTATUS,
    PHYEMAC0RXCHARISCOMMA,
    PHYEMAC0RXCHARISK,
    PHYEMAC0RXCHECKINGCRC,
    PHYEMAC0RXCLK,
    PHYEMAC0RXCLKCORCNT,
    PHYEMAC0RXCOMMADET,
    PHYEMAC0RXD,
    PHYEMAC0RXDISPERR,
    PHYEMAC0RXDV,
    PHYEMAC0RXER,
    PHYEMAC0RXLOSSOFSYNC,
    PHYEMAC0RXNOTINTABLE,
    PHYEMAC0RXRUNDISP,
    PHYEMAC0SIGNALDET,
    PHYEMAC0TXBUFERR,
    PHYEMAC1COL,
    PHYEMAC1CRS,
    PHYEMAC1GTXCLK,
    PHYEMAC1MCLKIN,
    PHYEMAC1MDIN,
    PHYEMAC1MIITXCLK,
    PHYEMAC1PHYAD,
    PHYEMAC1RXBUFERR,
    PHYEMAC1RXBUFSTATUS,
    PHYEMAC1RXCHARISCOMMA,
    PHYEMAC1RXCHARISK,
    PHYEMAC1RXCHECKINGCRC,
    PHYEMAC1RXCLK,
    PHYEMAC1RXCLKCORCNT,
    PHYEMAC1RXCOMMADET,
    PHYEMAC1RXD,
    PHYEMAC1RXDISPERR,
    PHYEMAC1RXDV,
    PHYEMAC1RXER,
    PHYEMAC1RXLOSSOFSYNC,
    PHYEMAC1RXNOTINTABLE,
    PHYEMAC1RXRUNDISP,
    PHYEMAC1SIGNALDET,
    PHYEMAC1TXBUFERR,
    RESET,
    TIEEMAC0CONFIGVEC,
    TIEEMAC0UNICASTADDR,
    TIEEMAC1CONFIGVEC,
    TIEEMAC1UNICASTADDR
);
parameter LOC = "UNPLACED";
parameter EMAC0_MODE = "RGMII";
parameter EMAC1_MODE = "RGMII";
output DCRHOSTDONEIR;
output EMAC0CLIENTANINTERRUPT;
output EMAC0CLIENTRXBADFRAME;
output EMAC0CLIENTRXCLIENTCLKOUT;
output EMAC0CLIENTRXDVLD;
output EMAC0CLIENTRXDVLDMSW;
output EMAC0CLIENTRXDVREG6;
output EMAC0CLIENTRXFRAMEDROP;
output EMAC0CLIENTRXGOODFRAME;
output EMAC0CLIENTRXSTATSBYTEVLD;
output EMAC0CLIENTRXSTATSVLD;
output EMAC0CLIENTTXACK;
output EMAC0CLIENTTXCLIENTCLKOUT;
output EMAC0CLIENTTXCOLLISION;
output EMAC0CLIENTTXGMIIMIICLKOUT;
output EMAC0CLIENTTXRETRANSMIT;
output EMAC0CLIENTTXSTATS;
output EMAC0CLIENTTXSTATSBYTEVLD;
output EMAC0CLIENTTXSTATSVLD;
output EMAC0PHYENCOMMAALIGN;
output EMAC0PHYLOOPBACKMSB;
output EMAC0PHYMCLKOUT;
output EMAC0PHYMDOUT;
output EMAC0PHYMDTRI;
output EMAC0PHYMGTRXRESET;
output EMAC0PHYMGTTXRESET;
output EMAC0PHYPOWERDOWN;
output EMAC0PHYSYNCACQSTATUS;
output EMAC0PHYTXCHARDISPMODE;
output EMAC0PHYTXCHARDISPVAL;
output EMAC0PHYTXCHARISK;
output EMAC0PHYTXCLK;
output EMAC0PHYTXEN;
output EMAC0PHYTXER;
output EMAC1CLIENTANINTERRUPT;
output EMAC1CLIENTRXBADFRAME;
output EMAC1CLIENTRXCLIENTCLKOUT;
output EMAC1CLIENTRXDVLD;
output EMAC1CLIENTRXDVLDMSW;
output EMAC1CLIENTRXDVREG6;
output EMAC1CLIENTRXFRAMEDROP;
output EMAC1CLIENTRXGOODFRAME;
output EMAC1CLIENTRXSTATSBYTEVLD;
output EMAC1CLIENTRXSTATSVLD;
output EMAC1CLIENTTXACK;
output EMAC1CLIENTTXCLIENTCLKOUT;
output EMAC1CLIENTTXCOLLISION;
output EMAC1CLIENTTXGMIIMIICLKOUT;
output EMAC1CLIENTTXRETRANSMIT;
output EMAC1CLIENTTXSTATS;
output EMAC1CLIENTTXSTATSBYTEVLD;
output EMAC1CLIENTTXSTATSVLD;
output EMAC1PHYENCOMMAALIGN;
output EMAC1PHYLOOPBACKMSB;
output EMAC1PHYMCLKOUT;
output EMAC1PHYMDOUT;
output EMAC1PHYMDTRI;
output EMAC1PHYMGTRXRESET;
output EMAC1PHYMGTTXRESET;
output EMAC1PHYPOWERDOWN;
output EMAC1PHYSYNCACQSTATUS;
output EMAC1PHYTXCHARDISPMODE;
output EMAC1PHYTXCHARDISPVAL;
output EMAC1PHYTXCHARISK;
output EMAC1PHYTXCLK;
output EMAC1PHYTXEN;
output EMAC1PHYTXER;
output EMACDCRACK;
output HOSTMIIMRDY;
output [0:31] EMACDCRDBUS;
output [15:0] EMAC0CLIENTRXD;
output [15:0] EMAC1CLIENTRXD;
output [31:0] HOSTRDDATA;
output [6:0] EMAC0CLIENTRXSTATS;
output [6:0] EMAC1CLIENTRXSTATS;
output [7:0] EMAC0PHYTXD;
output [7:0] EMAC1PHYTXD;
input CLIENTEMAC0DCMLOCKED;
input CLIENTEMAC0PAUSEREQ;
input CLIENTEMAC0RXCLIENTCLKIN;
input CLIENTEMAC0TXCLIENTCLKIN;
input CLIENTEMAC0TXDVLD;
input CLIENTEMAC0TXDVLDMSW;
input CLIENTEMAC0TXFIRSTBYTE;
input CLIENTEMAC0TXGMIIMIICLKIN;
input CLIENTEMAC0TXUNDERRUN;
input CLIENTEMAC1DCMLOCKED;
input CLIENTEMAC1PAUSEREQ;
input CLIENTEMAC1RXCLIENTCLKIN;
input CLIENTEMAC1TXCLIENTCLKIN;
input CLIENTEMAC1TXDVLD;
input CLIENTEMAC1TXDVLDMSW;
input CLIENTEMAC1TXFIRSTBYTE;
input CLIENTEMAC1TXGMIIMIICLKIN;
input CLIENTEMAC1TXUNDERRUN;
input DCREMACCLK;
input DCREMACENABLE;
input DCREMACREAD;
input DCREMACWRITE;
input HOSTCLK;
input HOSTEMAC1SEL;
input HOSTMIIMSEL;
input HOSTREQ;
input PHYEMAC0COL;
input PHYEMAC0CRS;
input PHYEMAC0GTXCLK;
input PHYEMAC0MCLKIN;
input PHYEMAC0MDIN;
input PHYEMAC0MIITXCLK;
input PHYEMAC0RXBUFERR;
input PHYEMAC0RXCHARISCOMMA;
input PHYEMAC0RXCHARISK;
input PHYEMAC0RXCHECKINGCRC;
input PHYEMAC0RXCLK;
input PHYEMAC0RXCOMMADET;
input PHYEMAC0RXDISPERR;
input PHYEMAC0RXDV;
input PHYEMAC0RXER;
input PHYEMAC0RXNOTINTABLE;
input PHYEMAC0RXRUNDISP;
input PHYEMAC0SIGNALDET;
input PHYEMAC0TXBUFERR;
input PHYEMAC1COL;
input PHYEMAC1CRS;
input PHYEMAC1GTXCLK;
input PHYEMAC1MCLKIN;
input PHYEMAC1MDIN;
input PHYEMAC1MIITXCLK;
input PHYEMAC1RXBUFERR;
input PHYEMAC1RXCHARISCOMMA;
input PHYEMAC1RXCHARISK;
input PHYEMAC1RXCHECKINGCRC;
input PHYEMAC1RXCLK;
input PHYEMAC1RXCOMMADET;
input PHYEMAC1RXDISPERR;
input PHYEMAC1RXDV;
input PHYEMAC1RXER;
input PHYEMAC1RXNOTINTABLE;
input PHYEMAC1RXRUNDISP;
input PHYEMAC1SIGNALDET;
input PHYEMAC1TXBUFERR;
input RESET;
input [0:31] DCREMACDBUS;
input [15:0] CLIENTEMAC0PAUSEVAL;
input [15:0] CLIENTEMAC0TXD;
input [15:0] CLIENTEMAC1PAUSEVAL;
input [15:0] CLIENTEMAC1TXD;
input [1:0] HOSTOPCODE;
input [1:0] PHYEMAC0RXBUFSTATUS;
input [1:0] PHYEMAC0RXLOSSOFSYNC;
input [1:0] PHYEMAC1RXBUFSTATUS;
input [1:0] PHYEMAC1RXLOSSOFSYNC;
input [2:0] PHYEMAC0RXCLKCORCNT;
input [2:0] PHYEMAC1RXCLKCORCNT;
input [31:0] HOSTWRDATA;
input [47:0] TIEEMAC0UNICASTADDR;
input [47:0] TIEEMAC1UNICASTADDR;
input [4:0] PHYEMAC0PHYAD;
input [4:0] PHYEMAC1PHYAD;
input [79:0] TIEEMAC0CONFIGVEC;
input [79:0] TIEEMAC1CONFIGVEC;
input [7:0] CLIENTEMAC0TXIFGDELAY;
input [7:0] CLIENTEMAC1TXIFGDELAY;
input [7:0] PHYEMAC0RXD;
input [7:0] PHYEMAC1RXD;
input [8:9] DCREMACABUS;
input [9:0] HOSTADDR;

endmodule
