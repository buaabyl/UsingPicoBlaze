// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/xec_libs/data/unisims/PPC440.v,v 1.2 2007/12/07 01:01:21 vandanad Exp $
///////////////////////////////////////////////////////////
//  Copyright (c) 1995/2006 Xilinx Inc.
//  All Right Reserved.
///////////////////////////////////////////////////////////
//
//   ____   ___
//  /   /\/   / 
// /___/  \  /    Vendor      : Xilinx 
// \  \    \/     Version : 10.1
//  \  \          Description : 
//  /  /                      
// /__/   /\      Filename    : PPC440.v
// \  \  /  \     Timestamp   : Thu Apr 19 10:07:12 2007

//  \__\/\__ \                    
//                                 
///////////////////////////////////////////////////////////

`timescale 1 ps / 1 ps 

module PPC440 (
    APUFCMDECFPUOP,
    APUFCMDECLDSTXFERSIZE,
    APUFCMDECLOAD,
    APUFCMDECNONAUTON,
    APUFCMDECSTORE,
    APUFCMDECUDI,
    APUFCMDECUDIVALID,
    APUFCMENDIAN,
    APUFCMFLUSH,
    APUFCMINSTRUCTION,
    APUFCMINSTRVALID,
    APUFCMLOADBYTEADDR,
    APUFCMLOADDATA,
    APUFCMLOADDVALID,
    APUFCMMSRFE0,
    APUFCMMSRFE1,
    APUFCMNEXTINSTRREADY,
    APUFCMOPERANDVALID,
    APUFCMRADATA,
    APUFCMRBDATA,
    APUFCMWRITEBACKOK,
    C440CPMCORESLEEPREQ,
    C440CPMDECIRPTREQ,
    C440CPMFITIRPTREQ,
    C440CPMMSRCE,
    C440CPMMSREE,
    C440CPMTIMERRESETREQ,
    C440CPMWDIRPTREQ,
    C440DBGSYSTEMCONTROL,
    C440JTGTDO,
    C440JTGTDOEN,
    C440MACHINECHECK,
    C440RSTCHIPRESETREQ,
    C440RSTCORERESETREQ,
    C440RSTSYSTEMRESETREQ,
    C440TRCBRANCHSTATUS,
    C440TRCCYCLE,
    C440TRCEXECUTIONSTATUS,
    C440TRCTRACESTATUS,
    C440TRCTRIGGEREVENTOUT,
    C440TRCTRIGGEREVENTTYPE,
    DMA0LLRSTENGINEACK,
    DMA0LLRXDSTRDYN,
    DMA0LLTXD,
    DMA0LLTXEOFN,
    DMA0LLTXEOPN,
    DMA0LLTXREM,
    DMA0LLTXSOFN,
    DMA0LLTXSOPN,
    DMA0LLTXSRCRDYN,
    DMA0RXIRQ,
    DMA0TXIRQ,
    DMA1LLRSTENGINEACK,
    DMA1LLRXDSTRDYN,
    DMA1LLTXD,
    DMA1LLTXEOFN,
    DMA1LLTXEOPN,
    DMA1LLTXREM,
    DMA1LLTXSOFN,
    DMA1LLTXSOPN,
    DMA1LLTXSRCRDYN,
    DMA1RXIRQ,
    DMA1TXIRQ,
    DMA2LLRSTENGINEACK,
    DMA2LLRXDSTRDYN,
    DMA2LLTXD,
    DMA2LLTXEOFN,
    DMA2LLTXEOPN,
    DMA2LLTXREM,
    DMA2LLTXSOFN,
    DMA2LLTXSOPN,
    DMA2LLTXSRCRDYN,
    DMA2RXIRQ,
    DMA2TXIRQ,
    DMA3LLRSTENGINEACK,
    DMA3LLRXDSTRDYN,
    DMA3LLTXD,
    DMA3LLTXEOFN,
    DMA3LLTXEOPN,
    DMA3LLTXREM,
    DMA3LLTXSOFN,
    DMA3LLTXSOPN,
    DMA3LLTXSRCRDYN,
    DMA3RXIRQ,
    DMA3TXIRQ,
    MIMCADDRESS,
    MIMCADDRESSVALID,
    MIMCBANKCONFLICT,
    MIMCBYTEENABLE,
    MIMCREADNOTWRITE,
    MIMCROWCONFLICT,
    MIMCWRITEDATA,
    MIMCWRITEDATAVALID,
    PPCCPMINTERCONNECTBUSY,
    PPCDMDCRABUS,
    PPCDMDCRDBUSOUT,
    PPCDMDCRREAD,
    PPCDMDCRUABUS,
    PPCDMDCRWRITE,
    PPCDSDCRACK,
    PPCDSDCRDBUSIN,
    PPCDSDCRTIMEOUTWAIT,
    PPCEICINTERCONNECTIRQ,
    PPCMPLBABORT,
    PPCMPLBABUS,
    PPCMPLBBE,
    PPCMPLBBUSLOCK,
    PPCMPLBLOCKERR,
    PPCMPLBPRIORITY,
    PPCMPLBRDBURST,
    PPCMPLBREQUEST,
    PPCMPLBRNW,
    PPCMPLBSIZE,
    PPCMPLBTATTRIBUTE,
    PPCMPLBTYPE,
    PPCMPLBUABUS,
    PPCMPLBWRBURST,
    PPCMPLBWRDBUS,
    PPCS0PLBADDRACK,
    PPCS0PLBMBUSY,
    PPCS0PLBMIRQ,
    PPCS0PLBMRDERR,
    PPCS0PLBMWRERR,
    PPCS0PLBRDBTERM,
    PPCS0PLBRDCOMP,
    PPCS0PLBRDDACK,
    PPCS0PLBRDDBUS,
    PPCS0PLBRDWDADDR,
    PPCS0PLBREARBITRATE,
    PPCS0PLBSSIZE,
    PPCS0PLBWAIT,
    PPCS0PLBWRBTERM,
    PPCS0PLBWRCOMP,
    PPCS0PLBWRDACK,
    PPCS1PLBADDRACK,
    PPCS1PLBMBUSY,
    PPCS1PLBMIRQ,
    PPCS1PLBMRDERR,
    PPCS1PLBMWRERR,
    PPCS1PLBRDBTERM,
    PPCS1PLBRDCOMP,
    PPCS1PLBRDDACK,
    PPCS1PLBRDDBUS,
    PPCS1PLBRDWDADDR,
    PPCS1PLBREARBITRATE,
    PPCS1PLBSSIZE,
    PPCS1PLBWAIT,
    PPCS1PLBWRBTERM,
    PPCS1PLBWRCOMP,
    PPCS1PLBWRDACK,

    CPMC440CLK,
    CPMC440CLKEN,
    CPMC440CORECLOCKINACTIVE,
    CPMC440TIMERCLOCK,
    CPMDCRCLK,
    CPMDMA0LLCLK,
    CPMDMA1LLCLK,
    CPMDMA2LLCLK,
    CPMDMA3LLCLK,
    CPMFCMCLK,
    CPMINTERCONNECTCLK,
    CPMINTERCONNECTCLKEN,
    CPMINTERCONNECTCLKNTO1,
    CPMMCCLK,
    CPMPPCMPLBCLK,
    CPMPPCS0PLBCLK,
    CPMPPCS1PLBCLK,
    DBGC440DEBUGHALT,
    DBGC440SYSTEMSTATUS,
    DBGC440UNCONDDEBUGEVENT,
    DCRPPCDMACK,
    DCRPPCDMDBUSIN,
    DCRPPCDMTIMEOUTWAIT,
    DCRPPCDSABUS,
    DCRPPCDSDBUSOUT,
    DCRPPCDSREAD,
    DCRPPCDSWRITE,
    EICC440CRITIRQ,
    EICC440EXTIRQ,
    FCMAPUCONFIRMINSTR,
    FCMAPUCR,
    FCMAPUDONE,
    FCMAPUEXCEPTION,
    FCMAPUFPSCRFEX,
    FCMAPURESULT,
    FCMAPURESULTVALID,
    FCMAPUSLEEPNOTREADY,
    FCMAPUSTOREDATA,
    JTGC440TCK,
    JTGC440TDI,
    JTGC440TMS,
    JTGC440TRSTNEG,
    LLDMA0RSTENGINEREQ,
    LLDMA0RXD,
    LLDMA0RXEOFN,
    LLDMA0RXEOPN,
    LLDMA0RXREM,
    LLDMA0RXSOFN,
    LLDMA0RXSOPN,
    LLDMA0RXSRCRDYN,
    LLDMA0TXDSTRDYN,
    LLDMA1RSTENGINEREQ,
    LLDMA1RXD,
    LLDMA1RXEOFN,
    LLDMA1RXEOPN,
    LLDMA1RXREM,
    LLDMA1RXSOFN,
    LLDMA1RXSOPN,
    LLDMA1RXSRCRDYN,
    LLDMA1TXDSTRDYN,
    LLDMA2RSTENGINEREQ,
    LLDMA2RXD,
    LLDMA2RXEOFN,
    LLDMA2RXEOPN,
    LLDMA2RXREM,
    LLDMA2RXSOFN,
    LLDMA2RXSOPN,
    LLDMA2RXSRCRDYN,
    LLDMA2TXDSTRDYN,
    LLDMA3RSTENGINEREQ,
    LLDMA3RXD,
    LLDMA3RXEOFN,
    LLDMA3RXEOPN,
    LLDMA3RXREM,
    LLDMA3RXSOFN,
    LLDMA3RXSOPN,
    LLDMA3RXSRCRDYN,
    LLDMA3TXDSTRDYN,
    MCMIADDRREADYTOACCEPT,
    MCMIREADDATA,
    MCMIREADDATAERR,
    MCMIREADDATAVALID,
    PLBPPCMADDRACK,
    PLBPPCMMBUSY,
    PLBPPCMMIRQ,
    PLBPPCMMRDERR,
    PLBPPCMMWRERR,
    PLBPPCMRDBTERM,
    PLBPPCMRDDACK,
    PLBPPCMRDDBUS,
    PLBPPCMRDPENDPRI,
    PLBPPCMRDPENDREQ,
    PLBPPCMRDWDADDR,
    PLBPPCMREARBITRATE,
    PLBPPCMREQPRI,
    PLBPPCMSSIZE,
    PLBPPCMTIMEOUT,
    PLBPPCMWRBTERM,
    PLBPPCMWRDACK,
    PLBPPCMWRPENDPRI,
    PLBPPCMWRPENDREQ,
    PLBPPCS0ABORT,
    PLBPPCS0ABUS,
    PLBPPCS0BE,
    PLBPPCS0BUSLOCK,
    PLBPPCS0LOCKERR,
    PLBPPCS0MASTERID,
    PLBPPCS0MSIZE,
    PLBPPCS0PAVALID,
    PLBPPCS0RDBURST,
    PLBPPCS0RDPENDPRI,
    PLBPPCS0RDPENDREQ,
    PLBPPCS0RDPRIM,
    PLBPPCS0REQPRI,
    PLBPPCS0RNW,
    PLBPPCS0SAVALID,
    PLBPPCS0SIZE,
    PLBPPCS0TATTRIBUTE,
    PLBPPCS0TYPE,
    PLBPPCS0UABUS,
    PLBPPCS0WRBURST,
    PLBPPCS0WRDBUS,
    PLBPPCS0WRPENDPRI,
    PLBPPCS0WRPENDREQ,
    PLBPPCS0WRPRIM,
    PLBPPCS1ABORT,
    PLBPPCS1ABUS,
    PLBPPCS1BE,
    PLBPPCS1BUSLOCK,
    PLBPPCS1LOCKERR,
    PLBPPCS1MASTERID,
    PLBPPCS1MSIZE,
    PLBPPCS1PAVALID,
    PLBPPCS1RDBURST,
    PLBPPCS1RDPENDPRI,
    PLBPPCS1RDPENDREQ,
    PLBPPCS1RDPRIM,
    PLBPPCS1REQPRI,
    PLBPPCS1RNW,
    PLBPPCS1SAVALID,
    PLBPPCS1SIZE,
    PLBPPCS1TATTRIBUTE,
    PLBPPCS1TYPE,
    PLBPPCS1UABUS,
    PLBPPCS1WRBURST,
    PLBPPCS1WRDBUS,
    PLBPPCS1WRPENDPRI,
    PLBPPCS1WRPENDREQ,
    PLBPPCS1WRPRIM,
    RSTC440RESETCHIP,
    RSTC440RESETCORE,
    RSTC440RESETSYSTEM,
    TIEC440DCURDLDCACHEPLBPRIO,
    TIEC440DCURDNONCACHEPLBPRIO,
    TIEC440DCURDTOUCHPLBPRIO,
    TIEC440DCURDURGENTPLBPRIO,
    TIEC440DCUWRFLUSHPLBPRIO,
    TIEC440DCUWRSTOREPLBPRIO,
    TIEC440DCUWRURGENTPLBPRIO,
    TIEC440ENDIANRESET,
    TIEC440ERPNRESET,
    TIEC440ICURDFETCHPLBPRIO,
    TIEC440ICURDSPECPLBPRIO,
    TIEC440ICURDTOUCHPLBPRIO,
    TIEC440PIR,
    TIEC440PVR,
    TIEC440USERRESET,
    TIEDCRBASEADDR,
    TRCC440TRACEDISABLE,
    TRCC440TRIGGEREVENTIN

);

parameter CLOCK_DELAY = "FALSE";
parameter DCR_AUTOLOCK_ENABLE = "TRUE";
parameter PPCDM_ASYNCMODE = "FALSE";
parameter PPCDS_ASYNCMODE = "FALSE";
parameter PPCS0_WIDTH_128N64 = "TRUE";
parameter PPCS1_WIDTH_128N64 = "TRUE";
parameter [0:16] APU_CONTROL = 17'h02000;
parameter [0:23] APU_UDI0 = 24'h000000;
parameter [0:23] APU_UDI1 = 24'h000000;
parameter [0:23] APU_UDI10 = 24'h000000;
parameter [0:23] APU_UDI11 = 24'h000000;
parameter [0:23] APU_UDI12 = 24'h000000;
parameter [0:23] APU_UDI13 = 24'h000000;
parameter [0:23] APU_UDI14 = 24'h000000;
parameter [0:23] APU_UDI15 = 24'h000000;
parameter [0:23] APU_UDI2 = 24'h000000;
parameter [0:23] APU_UDI3 = 24'h000000;
parameter [0:23] APU_UDI4 = 24'h000000;
parameter [0:23] APU_UDI5 = 24'h000000;
parameter [0:23] APU_UDI6 = 24'h000000;
parameter [0:23] APU_UDI7 = 24'h000000;
parameter [0:23] APU_UDI8 = 24'h000000;
parameter [0:23] APU_UDI9 = 24'h000000;
parameter [0:31] DMA0_RXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA0_TXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA1_RXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA1_TXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA2_RXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA2_TXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA3_RXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA3_TXCHANNELCTRL = 32'h01010000;
parameter [0:31] INTERCONNECT_IMASK = 32'hFFFFFFFF;
parameter [0:31] INTERCONNECT_TMPL_SEL = 32'h3FFFFFFF;
parameter [0:31] MI_ARBCONFIG = 32'h00432010;
parameter [0:31] MI_BANKCONFLICT_MASK = 32'h00000000;
parameter [0:31] MI_CONTROL = 32'h0000008F;
parameter [0:31] MI_ROWCONFLICT_MASK = 32'h00000000;
parameter [0:31] PPCM_ARBCONFIG = 32'h00432010;
parameter [0:31] PPCM_CONTROL = 32'h8000019F;
parameter [0:31] PPCM_COUNTER = 32'h00000500;
parameter [0:31] PPCS0_ADDRMAP_TMPL0 = 32'hFFFFFFFF;
parameter [0:31] PPCS0_ADDRMAP_TMPL1 = 32'hFFFFFFFF;
parameter [0:31] PPCS0_ADDRMAP_TMPL2 = 32'hFFFFFFFF;
parameter [0:31] PPCS0_ADDRMAP_TMPL3 = 32'hFFFFFFFF;
parameter [0:31] PPCS0_CONTROL = 32'h8033336C;
parameter [0:31] PPCS1_ADDRMAP_TMPL0 = 32'hFFFFFFFF;
parameter [0:31] PPCS1_ADDRMAP_TMPL1 = 32'hFFFFFFFF;
parameter [0:31] PPCS1_ADDRMAP_TMPL2 = 32'hFFFFFFFF;
parameter [0:31] PPCS1_ADDRMAP_TMPL3 = 32'hFFFFFFFF;
parameter [0:31] PPCS1_CONTROL = 32'h8033336C;
parameter [0:31] XBAR_ADDRMAP_TMPL0 = 32'hFFFF0000;
parameter [0:31] XBAR_ADDRMAP_TMPL1 = 32'h00000000;
parameter [0:31] XBAR_ADDRMAP_TMPL2 = 32'h00000000;
parameter [0:31] XBAR_ADDRMAP_TMPL3 = 32'h00000000;
parameter [0:7] DMA0_CONTROL = 8'h00;
parameter [0:7] DMA1_CONTROL = 8'h00;
parameter [0:7] DMA2_CONTROL = 8'h00;
parameter [0:7] DMA3_CONTROL = 8'h00;
parameter [0:9] DMA0_RXIRQTIMER = 10'h3FF;
parameter [0:9] DMA0_TXIRQTIMER = 10'h3FF;
parameter [0:9] DMA1_RXIRQTIMER = 10'h3FF;
parameter [0:9] DMA1_TXIRQTIMER = 10'h3FF;
parameter [0:9] DMA2_RXIRQTIMER = 10'h3FF;
parameter [0:9] DMA2_TXIRQTIMER = 10'h3FF;
parameter [0:9] DMA3_RXIRQTIMER = 10'h3FF;
parameter [0:9] DMA3_TXIRQTIMER = 10'h3FF;

output APUFCMDECFPUOP;
output APUFCMDECLOAD;
output APUFCMDECNONAUTON;
output APUFCMDECSTORE;
output APUFCMDECUDIVALID;
output APUFCMENDIAN;
output APUFCMFLUSH;
output APUFCMINSTRVALID;
output APUFCMLOADDVALID;
output APUFCMMSRFE0;
output APUFCMMSRFE1;
output APUFCMNEXTINSTRREADY;
output APUFCMOPERANDVALID;
output APUFCMWRITEBACKOK;
output C440CPMCORESLEEPREQ;
output C440CPMDECIRPTREQ;
output C440CPMFITIRPTREQ;
output C440CPMMSRCE;
output C440CPMMSREE;
output C440CPMTIMERRESETREQ;
output C440CPMWDIRPTREQ;
output C440JTGTDO;
output C440JTGTDOEN;
output C440MACHINECHECK;
output C440RSTCHIPRESETREQ;
output C440RSTCORERESETREQ;
output C440RSTSYSTEMRESETREQ;
output C440TRCCYCLE;
output C440TRCTRIGGEREVENTOUT;
output DMA0LLRSTENGINEACK;
output DMA0LLRXDSTRDYN;
output DMA0LLTXEOFN;
output DMA0LLTXEOPN;
output DMA0LLTXSOFN;
output DMA0LLTXSOPN;
output DMA0LLTXSRCRDYN;
output DMA0RXIRQ;
output DMA0TXIRQ;
output DMA1LLRSTENGINEACK;
output DMA1LLRXDSTRDYN;
output DMA1LLTXEOFN;
output DMA1LLTXEOPN;
output DMA1LLTXSOFN;
output DMA1LLTXSOPN;
output DMA1LLTXSRCRDYN;
output DMA1RXIRQ;
output DMA1TXIRQ;
output DMA2LLRSTENGINEACK;
output DMA2LLRXDSTRDYN;
output DMA2LLTXEOFN;
output DMA2LLTXEOPN;
output DMA2LLTXSOFN;
output DMA2LLTXSOPN;
output DMA2LLTXSRCRDYN;
output DMA2RXIRQ;
output DMA2TXIRQ;
output DMA3LLRSTENGINEACK;
output DMA3LLRXDSTRDYN;
output DMA3LLTXEOFN;
output DMA3LLTXEOPN;
output DMA3LLTXSOFN;
output DMA3LLTXSOPN;
output DMA3LLTXSRCRDYN;
output DMA3RXIRQ;
output DMA3TXIRQ;
output MIMCADDRESSVALID;
output MIMCBANKCONFLICT;
output MIMCREADNOTWRITE;
output MIMCROWCONFLICT;
output MIMCWRITEDATAVALID;
output PPCCPMINTERCONNECTBUSY;
output PPCDMDCRREAD;
output PPCDMDCRWRITE;
output PPCDSDCRACK;
output PPCDSDCRTIMEOUTWAIT;
output PPCEICINTERCONNECTIRQ;
output PPCMPLBABORT;
output PPCMPLBBUSLOCK;
output PPCMPLBLOCKERR;
output PPCMPLBRDBURST;
output PPCMPLBREQUEST;
output PPCMPLBRNW;
output PPCMPLBWRBURST;
output PPCS0PLBADDRACK;
output PPCS0PLBRDBTERM;
output PPCS0PLBRDCOMP;
output PPCS0PLBRDDACK;
output PPCS0PLBREARBITRATE;
output PPCS0PLBWAIT;
output PPCS0PLBWRBTERM;
output PPCS0PLBWRCOMP;
output PPCS0PLBWRDACK;
output PPCS1PLBADDRACK;
output PPCS1PLBRDBTERM;
output PPCS1PLBRDCOMP;
output PPCS1PLBRDDACK;
output PPCS1PLBREARBITRATE;
output PPCS1PLBWAIT;
output PPCS1PLBWRBTERM;
output PPCS1PLBWRCOMP;
output PPCS1PLBWRDACK;
output [0:127] APUFCMLOADDATA;
output [0:127] MIMCWRITEDATA;
output [0:127] PPCMPLBWRDBUS;
output [0:127] PPCS0PLBRDDBUS;
output [0:127] PPCS1PLBRDDBUS;
output [0:13] C440TRCTRIGGEREVENTTYPE;
output [0:15] MIMCBYTEENABLE;
output [0:15] PPCMPLBBE;
output [0:15] PPCMPLBTATTRIBUTE;
output [0:1] PPCMPLBPRIORITY;
output [0:1] PPCS0PLBSSIZE;
output [0:1] PPCS1PLBSSIZE;
output [0:2] APUFCMDECLDSTXFERSIZE;
output [0:2] C440TRCBRANCHSTATUS;
output [0:2] PPCMPLBTYPE;
output [0:31] APUFCMINSTRUCTION;
output [0:31] APUFCMRADATA;
output [0:31] APUFCMRBDATA;
output [0:31] DMA0LLTXD;
output [0:31] DMA1LLTXD;
output [0:31] DMA2LLTXD;
output [0:31] DMA3LLTXD;
output [0:31] PPCDMDCRDBUSOUT;
output [0:31] PPCDSDCRDBUSIN;
output [0:31] PPCMPLBABUS;
output [0:35] MIMCADDRESS;
output [0:3] APUFCMDECUDI;
output [0:3] APUFCMLOADBYTEADDR;
output [0:3] DMA0LLTXREM;
output [0:3] DMA1LLTXREM;
output [0:3] DMA2LLTXREM;
output [0:3] DMA3LLTXREM;
output [0:3] PPCMPLBSIZE;
output [0:3] PPCS0PLBMBUSY;
output [0:3] PPCS0PLBMIRQ;
output [0:3] PPCS0PLBMRDERR;
output [0:3] PPCS0PLBMWRERR;
output [0:3] PPCS0PLBRDWDADDR;
output [0:3] PPCS1PLBMBUSY;
output [0:3] PPCS1PLBMIRQ;
output [0:3] PPCS1PLBMRDERR;
output [0:3] PPCS1PLBMWRERR;
output [0:3] PPCS1PLBRDWDADDR;
output [0:4] C440TRCEXECUTIONSTATUS;
output [0:6] C440TRCTRACESTATUS;
output [0:7] C440DBGSYSTEMCONTROL;
output [0:9] PPCDMDCRABUS;
output [20:21] PPCDMDCRUABUS;
output [28:31] PPCMPLBUABUS;

input CPMC440CLK;
input CPMC440CLKEN;
input CPMC440CORECLOCKINACTIVE;
input CPMC440TIMERCLOCK;
input CPMDCRCLK;
input CPMDMA0LLCLK;
input CPMDMA1LLCLK;
input CPMDMA2LLCLK;
input CPMDMA3LLCLK;
input CPMFCMCLK;
input CPMINTERCONNECTCLK;
input CPMINTERCONNECTCLKEN;
input CPMINTERCONNECTCLKNTO1;
input CPMMCCLK;
input CPMPPCMPLBCLK;
input CPMPPCS0PLBCLK;
input CPMPPCS1PLBCLK;
input DBGC440DEBUGHALT;
input DBGC440UNCONDDEBUGEVENT;
input DCRPPCDMACK;
input DCRPPCDMTIMEOUTWAIT;
input DCRPPCDSREAD;
input DCRPPCDSWRITE;
input EICC440CRITIRQ;
input EICC440EXTIRQ;
input FCMAPUCONFIRMINSTR;
input FCMAPUDONE;
input FCMAPUEXCEPTION;
input FCMAPUFPSCRFEX;
input FCMAPURESULTVALID;
input FCMAPUSLEEPNOTREADY;
input JTGC440TCK;
input JTGC440TDI;
input JTGC440TMS;
input JTGC440TRSTNEG;
input LLDMA0RSTENGINEREQ;
input LLDMA0RXEOFN;
input LLDMA0RXEOPN;
input LLDMA0RXSOFN;
input LLDMA0RXSOPN;
input LLDMA0RXSRCRDYN;
input LLDMA0TXDSTRDYN;
input LLDMA1RSTENGINEREQ;
input LLDMA1RXEOFN;
input LLDMA1RXEOPN;
input LLDMA1RXSOFN;
input LLDMA1RXSOPN;
input LLDMA1RXSRCRDYN;
input LLDMA1TXDSTRDYN;
input LLDMA2RSTENGINEREQ;
input LLDMA2RXEOFN;
input LLDMA2RXEOPN;
input LLDMA2RXSOFN;
input LLDMA2RXSOPN;
input LLDMA2RXSRCRDYN;
input LLDMA2TXDSTRDYN;
input LLDMA3RSTENGINEREQ;
input LLDMA3RXEOFN;
input LLDMA3RXEOPN;
input LLDMA3RXSOFN;
input LLDMA3RXSOPN;
input LLDMA3RXSRCRDYN;
input LLDMA3TXDSTRDYN;
input MCMIADDRREADYTOACCEPT;
input MCMIREADDATAERR;
input MCMIREADDATAVALID;
input PLBPPCMADDRACK;
input PLBPPCMMBUSY;
input PLBPPCMMIRQ;
input PLBPPCMMRDERR;
input PLBPPCMMWRERR;
input PLBPPCMRDBTERM;
input PLBPPCMRDDACK;
input PLBPPCMRDPENDREQ;
input PLBPPCMREARBITRATE;
input PLBPPCMTIMEOUT;
input PLBPPCMWRBTERM;
input PLBPPCMWRDACK;
input PLBPPCMWRPENDREQ;
input PLBPPCS0ABORT;
input PLBPPCS0BUSLOCK;
input PLBPPCS0LOCKERR;
input PLBPPCS0PAVALID;
input PLBPPCS0RDBURST;
input PLBPPCS0RDPENDREQ;
input PLBPPCS0RDPRIM;
input PLBPPCS0RNW;
input PLBPPCS0SAVALID;
input PLBPPCS0WRBURST;
input PLBPPCS0WRPENDREQ;
input PLBPPCS0WRPRIM;
input PLBPPCS1ABORT;
input PLBPPCS1BUSLOCK;
input PLBPPCS1LOCKERR;
input PLBPPCS1PAVALID;
input PLBPPCS1RDBURST;
input PLBPPCS1RDPENDREQ;
input PLBPPCS1RDPRIM;
input PLBPPCS1RNW;
input PLBPPCS1SAVALID;
input PLBPPCS1WRBURST;
input PLBPPCS1WRPENDREQ;
input PLBPPCS1WRPRIM;
input RSTC440RESETCHIP;
input RSTC440RESETCORE;
input RSTC440RESETSYSTEM;
input TIEC440ENDIANRESET;
input TRCC440TRACEDISABLE;
input TRCC440TRIGGEREVENTIN;
input [0:127] FCMAPUSTOREDATA;
input [0:127] MCMIREADDATA;
input [0:127] PLBPPCMRDDBUS;
input [0:127] PLBPPCS0WRDBUS;
input [0:127] PLBPPCS1WRDBUS;
input [0:15] PLBPPCS0BE;
input [0:15] PLBPPCS0TATTRIBUTE;
input [0:15] PLBPPCS1BE;
input [0:15] PLBPPCS1TATTRIBUTE;
input [0:1] PLBPPCMRDPENDPRI;
input [0:1] PLBPPCMREQPRI;
input [0:1] PLBPPCMSSIZE;
input [0:1] PLBPPCMWRPENDPRI;
input [0:1] PLBPPCS0MASTERID;
input [0:1] PLBPPCS0MSIZE;
input [0:1] PLBPPCS0RDPENDPRI;
input [0:1] PLBPPCS0REQPRI;
input [0:1] PLBPPCS0WRPENDPRI;
input [0:1] PLBPPCS1MASTERID;
input [0:1] PLBPPCS1MSIZE;
input [0:1] PLBPPCS1RDPENDPRI;
input [0:1] PLBPPCS1REQPRI;
input [0:1] PLBPPCS1WRPENDPRI;
input [0:1] TIEC440DCURDLDCACHEPLBPRIO;
input [0:1] TIEC440DCURDNONCACHEPLBPRIO;
input [0:1] TIEC440DCURDTOUCHPLBPRIO;
input [0:1] TIEC440DCURDURGENTPLBPRIO;
input [0:1] TIEC440DCUWRFLUSHPLBPRIO;
input [0:1] TIEC440DCUWRSTOREPLBPRIO;
input [0:1] TIEC440DCUWRURGENTPLBPRIO;
input [0:1] TIEC440ICURDFETCHPLBPRIO;
input [0:1] TIEC440ICURDSPECPLBPRIO;
input [0:1] TIEC440ICURDTOUCHPLBPRIO;
input [0:1] TIEDCRBASEADDR;
input [0:2] PLBPPCS0TYPE;
input [0:2] PLBPPCS1TYPE;
input [0:31] DCRPPCDMDBUSIN;
input [0:31] DCRPPCDSDBUSOUT;
input [0:31] FCMAPURESULT;
input [0:31] LLDMA0RXD;
input [0:31] LLDMA1RXD;
input [0:31] LLDMA2RXD;
input [0:31] LLDMA3RXD;
input [0:31] PLBPPCS0ABUS;
input [0:31] PLBPPCS1ABUS;
input [0:3] FCMAPUCR;
input [0:3] LLDMA0RXREM;
input [0:3] LLDMA1RXREM;
input [0:3] LLDMA2RXREM;
input [0:3] LLDMA3RXREM;
input [0:3] PLBPPCMRDWDADDR;
input [0:3] PLBPPCS0SIZE;
input [0:3] PLBPPCS1SIZE;
input [0:3] TIEC440ERPNRESET;
input [0:3] TIEC440USERRESET;
input [0:4] DBGC440SYSTEMSTATUS;
input [0:9] DCRPPCDSABUS;
input [28:31] PLBPPCS0UABUS;
input [28:31] PLBPPCS1UABUS;
input [28:31] TIEC440PIR;
input [28:31] TIEC440PVR;

endmodule
